BZh91AY&SY���� �_�Pxg���������P�r](v�� �PzF��� �2   �4*~���4=L���1 � ��&M"�P��<(�h h���&L��L �0L�0�D�L���44&Q�?T� 4���R�hOzBH(�V$ ~?/3�"fq�hRi$א|(ۀ�hЬb�
%�n �a7{����6��+�L�,�RQ#�j�����֛�ڢ�$�29�:����|٧*l���0���FT�bA���^C+�"���yf�f[I�T=K����F�g���U:�^y�X���,�^͡��p^1"۰XהsX0�=R�|B�z>�eI���f%/�eU�"��f\l��-D��)A����7�C��KLfv�[J�\��(Rש�A�
<��9�H�[��J�f�Q�3u��XHBBΒI(��5��p�4�ߑˑ�%Q.Z�J(�Cu���Q��8���"0�����H j6���@$E�.q��z���1�������ᣏX��<`��iH�6�<��.�����.FI)s��W%�5�������xÐ;w.�����~a�FN���A�e;3��i�1L<����7e\��3&ԗ�iQX��r�y�`X&m`l^V$LcP�e��� �,̒xP%Zٓ9\�57h�A���I�ѹ�(�1i(9DL�)XR�qg5r���.����18�S~��`2�c� 񦥬4���XN�i���WN����!�A���$�Z���|&���T4RSB���bQl��$�Pe޷�l�fMZ/5���ֶ�̽5�Q��R{v↋��]�q�=�4s�[a��q�3�XKpT``L/h��V�4�^��f`0��φA!A�
�����%D��)��s*M�S�&TDM�q�n�܄��PF�`3���#�\lv&`�<	�����F�*��
@���\����&T<3�L�Q�Z���P�(6��3~�J��!���#n*3Vʆ�²dź��u�,'P����B�T�C �i3.%�jH6�9)m֒
X0�3��xUA��R�i�z�s�L\H9�����a�\U���q���F�;2,�4�
���nJ��H�
��8`