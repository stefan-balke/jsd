BZh91AY&SY�÷� _�Px���������P㵀r†5S�=M���H@4h2  �MS��P     hBDF�h6������  @0`��`ѐ��&��D��0D�	����=G��@(�<���OrB!	 
� ~>_��\� ��R`�!���_vZ7�`cB�34r�TH�Hg6j4�n������&v6d㢙D��|�޼o!X�u*�0��ێ����H��Jڀ�ABt��0 ,��p��%�|ٔ�'D\�v��f���T
��6��� �/��P`@��@����?��4ŃI��\̣
T�uK��ʕm)�0�3dh���`ނ4/
��O2��2���ܼ+%{�tq4��v*�&�!e�kc���tX�aJ���YQ{�؋�R����,0�o+[<�]LE��P���7v�m��B�ѯ�
KodC���*Q%�ڤx��1�q�P��6���d�n�8�C*�gD-�#[�YA�6H�U��1b:���ne� �0.~=W	T`��AT��{'���t���q�0@e3n,�
o�����H�:��%�@+��g�1`� 0���j�P���A|���[Q�*�FWjK��P�G�1� �y�(&m`k^U	��Ȱ;��>enI;�	R��f ��q��o��ȋ�Ţp5t2��L��P�"�ֈ���B;��KP�g�AR�������Ç df
���Aٟ�kFsJ�W�
��v���Y�R`�sH2$����tS ͖�dƺ����'��k�QH0S;������l���i��#�E�&(�zd�M)N;�#��`�i"T�#��� ��S�>�Ò��t�8%�(00&�Nf��7<g(��i @H�ҠE�;�,HHF/Q.�p�*C�3�2��Ҁ�l��f&�rʜ�:��fӀ�G���� ��Y�v�c�CBe9�a�*I!�9��w^�����b��<N������P�,NhÁ"�8D�K�~��Tf[7�*B)ho�`o����T,Sz-�X"���V����Ł��6|Ă�:K%�rT@��Ťa��`ki4�::N@�����ƵiQi� ݾ���6�M�u���H�d0hL�@srE8P��÷�