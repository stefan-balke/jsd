BZh91AY&SY�p �߀Px����������P��u�I��&AL%h�j4�)�2�@4h�� �I�Q� �  h    ��$�mL��h  @��b�LFCC �#I S#�iOd��=4ȍ14� �bq��+|D��a"2�K!^�w䫜���0bJ��F�ۘq�~l 3K ��j�$�d��{�����Ow�����ޭA��e��p���,�I�+r�6�Z��Tŉ�TMNa�à["4�y�H(�R୭��a[k��p�Ksm ����F@�)[�#��M%�Z�Y��3�GLG.G& AQAE����;n��Ų�%-:w����K�j������h�&&6��{&���Q+L2�-��T�\�yRf	�h���M�3<+�P2Z��P�.�k
pB�!T(
;@G*��`Gq��\wδ���Z���["�Y-U���y�:.���oB"�ɦ2��M\V�+`����b�
Jݦ"���	�v�Br�p��=��.y��<C8$1���m������m�rw�B�;�:%J$����C�dJr����(�j�6X�"F<a-�$vY���t-�PP0�u����Ũ��M�}ɖ>!�6�'@iO>�O�$�)������E!��Y)����a>�LH�QI*�{ޑYP��袥���Lܱ��ß�w{��þF���-J28�:��z��6�&�Ȳ�\?��ҋ�uOz���<s
���G�6Ss߁����sOu�(��6�|r=^ZYg���I[0.�t��F�o+��K9�h��7o��)��|��WXC���1�fb�ٿ�ևsp���uAР�f�V�#�zF���s��%�c�G����l�d�\X��,)K�j��u�c�"W9"B��q�aXQ�8� )7�ʂ}C���A�*�0��~�	��������-=�z;�⣃�v��9����5��t#k�U"�٘ڪ��֥�H
6�Ab��tHF��%�.�`Ρhnԭ�qSF�1%����`��[p�#��^)��$��|�ؾ�G�S�rE�O���#��u�%;�O�%��AJ:^M�k;#��k��8�]�&��Չ�Q�U+S~�.R��V�֋����^���p^�?FZ�F:NF��d[ ����R��(d#6�a�j
��.g���d�u�a�~�w��/f��ze��#?�q�n�(���ncECr.d�}4��v$[[-�UL����P*�API�?�]��B@Tz��