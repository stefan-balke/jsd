BZh91AY&SY�D,� n߀@x����������Px�6\�M� J!2��S���h4@ �F�SB4MP� �d i�   �����#F2	��3S ё�@�44�0&&�	�&L�&	����MM�d&MS�Ԟ����mF�����ʐ��i$���=_���Ȁ���*J���O͛pZ�$���D4gj�2D#	��7vv77|7<�3����Ρ9����Ԣ�-�y�	)"�tH�⃏�Y����וr�A�$`9R� Z�F�ĄI�<[�Mi�����Bj씐�@�^�d�@���J�����ǭW �1���N�Í�E~!m�Zl�A����V�ZB'�������6��3�W+���mĘk�AșԂ�����3.�I�˶V-�D��XO`{�3��5�j�E��A&5i5v�$��bd��&cTAQ�k�F���� �\�';a�kQ,E��f1*1f!b�$��.Q�����:gl\���!���oY��hhC�co@oP��#�
�=TJ�I.�X��mjwTnH��������vQ9uUQ@��a�Tt�[0@@ t�6�1�d&Hm}֡/��1~C����,����gW�3�o��h�/u4�s�и}\���#^/�I*���J�r�k����;D0�ǅ�g@3/�:����1q� ���&I��*�G 8�� :�	�)�䗥@u ��ɘ���@bf�k�T)"�|hg��?�Ή'|�4��'��Nz���Bg+c���dŹ4�X���a;��I�3�.C�χ"�oH!�1'D��¡K����h���A���#��>��,T�q�362K�"�G*dn=d���c$,�N�f�p`��d� ���K1
NE�d�T����DY��$���|���l �: ���x�0SP�����Ԩ0.$CA)
A�_'�\I$�3l�"��ج:$#A�K�,]�Je�冄���P��p};qG��'���s7�@2�J�����ˌ��\��Ǭ�x�b����|�!�2�O��"�}�`�E���6�bG�iS��X3�;�.
�4�dF4�NB�����Lf{w�*A��E��ĩ*�^�x �lH������PZ�L7Ю��
�`snq���J�IH����a�{03LG�@�Ȱ44��j҈/� n��n�m{ͪu���0c�n���]��BB��