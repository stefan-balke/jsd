BZh91AY&SY��0 �_�Py���������P�ꋱ�sR� D����=&�z�6S�z�� �?T�S�P�4     ���b=OSC��hhz� �̐q�&LF& L�&@F �"��d&������zCM 1D�f�C�@I@@'��s��T�n�26Ҕ�T�_�{E),E�M9aI0w1e%{�c�@��������gB�'4�̨c�Xf�ۭS��������KW,rG���r)����k���-)	 �u�Ԯ[����M��-�:F辽���T�i���M)z�J8c�M	L�pAo"؈h�M�%�<�%�_�M�d��\��0�Z�b4ڥ���ʈ���/*N�J�\ଋ�_A�TH � @-%m6-K3p��%$���4�+\�8Ʈ��u�46���V�i��ƹu>냏T;E"�k(9)��ô���s��ْ4�^	JC�D�L!����]�3�Ę���/鶿!�.�vհ�V�:�:n�O�BȱǙ�R������{���{ϓ��Tks%�i���of�&�Ds�#���ԙ�����O����bd���[o)wa֫:i,��O�`3�[Fg��F%�K�Hp9�P�*��ғ��(��V�W��tb��k�_v��ၖ��lK��7�Y����<�)nJi�P�n�9�4.*h҉s��P�%�{ʎ33a��̢�T��8����F���?r�Y��0�tA-g�9^e%�i*2��,��1���Ƭ$`�{O��f��1�0`^�
�F r�Ƣ����h�Ԭp��қ"a�A�w��C�4����-B�o���T��
:DCA튁Uj��bgZ��F�;(����4s⁩@7����d���i�&�Fy���x�|���P{���df�[��}�!��<�
�d�i��q�ä�o�4]5e6�f~.T���)>+�܍�x�] ��HƲ��
l�����M��岤����4�9(g��i���,YB�6�t�`hZ��fz��v<D\�`ms�`:��H�]�_<����[��y�����O����)��!��