BZh91AY&SY� í �_�Px���������`<u� չ�� p�JO�=��L��4A��A����Q@��=C126����&L�20�&�db``��*z	�Dh��{TS@  � 0&&�	�&L�&	�����$���L��4S��M��  �MO)��Es�-"I��4�E�����Uv�G��΢^*)z�'ኪ�|p��0F&L����%�f"#	�����,wI|&�k�N��G)�)���l��Oۓ��6�F� -�m��+��6z�	�"DEB��Q���aq���m%�\��S���I��5D�"(�v�1Ы�� ��"Hg�nI&f�ȝr�KEF���ſ|DU$/�X������,���;������?mӞ�<t�qߤ��!$��72-��5����Ú0C���0i�kƚ`v�����	7*D�l�7�u@�,�k3� ���ERU-ҭz.��ow��Kl;@J*K��>6-X��LE٨��(&L�f��!\���*��)w���3��G,h|�ξ��ʾ3����Ocb�4d�5�$�	ĭ2ښDS�"H�Z�,��\�b�1F���W�����*�������6��wTUm��Y,��;Rl�3=��Fs�b�PHB���U��I9�GWxw�#Ÿ�h��O���∪,��P$�D}%�^b!%	$`DDDK`�zJ��Je{�f5\�r�T�8���
��M̄�Y=+�q���(��@i�y���IFةS�h�O�����pO�~hjD�z9�����2�j�Օ��&U�6���F,XE��F�~�g������=���!�KB��c�^n��i�̥��q�Ϯ�8xO�O�W9'��DG�!�q|�2Jr��|�bT�Z�����K,����+�"�禭ќ1
�H#��b�1'L+-������|���S]�������=Y슲�/�L��TT�U��>��j��ގé��|�.f�������|��w����'vq������Ʌ��Q���{�v��N��d����m����n��q��C�l�R,[c�_Kտ<����*6Κ�u�̇���*=L�B�ڣ�F���~�9I4P���Rè��Xߋ�[aab���d\��Vy�q�0{�b�!Eˊ��1j�6ib�V���<yD�u��;�`S��t�R>�����.-�����w(�1;doj½�Z�S?���x�}�r(���Cy�0�o�/kQ���y�L�R�
ww)u(�U�����o+sjS��M���=�=q6��v�fb^�5�2!�]�Yk:�f�b����瑫�R�)[+�M�u�F#}�7)�uH�����5%���v8�v�8��rW�9s�04u�U7Ѯ�]!�P��G7�]��BB4�