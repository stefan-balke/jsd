BZh91AY&SY�ڬ� �߀Px���������P~p��+@VH�$�6��   h h4LL���       �)�=G�Hm@z���@�=@���&L�20�&�db``
�M�OM
yOSj6P� �M4ɱy"��KD�4D�B���`��TLB�T�aU^��5*&�̰�h�j�H$f@���:�n���ϋ�;{|���͗�1je˫��v��-]h��چ;��os�n�W��������(��m�5І��+�6�y���Щ�~V[�F����l �r�R��:g��{��L���m�.D0cׇ��<|"5\������8]bօ�����ze��[J�ջ'"j^D�h�h��a���@Wf�����{���"�8��:��1J����2jZ� !�́ ���0�L��h�fD��@�D)���/a[T-�)K��"���h*�	t�w(wB��A݄�I��֩E	��c�X���7���hi!��������#�B�;ϋ6*���u��z�XSc(`���V �2b���hA����A�P5�B��A@�5��|�4�aS����GS���!<ר�|��eG�_��Q�/S�dm�B��蘿�=!v��:�oT�TB4pp3M}9�{~�K�PU`NW$z�rA�Վ������$j�R�(X�mw׋n�2\�)hg���(,�_cZ�шP@q�4"��? :X^yH�c#9ˇ�{!#=�Jm�Vs���z4ǣ��y�숹]ܓ�j�S�GT��u��Mv�+L2[K���٧lU��v�5Mu[������h�W�n�F_'+R	�(�ge����6^�������/#N���o�*1��7ף3����]�S_�>��kN�\��uk�sR,X�����\!��C#I^d��B��3|F�������ݦ�F�FJ���/w)�����7@��Ab��$$#G޵�ȣQ�T�SB�vKŪ2<�k��-��rx�D�����t��3yf�#߇ˠ�spm,:���ৡ3y�W�r�%1�w8�HWP�Tv��~~n1����SC���v&�܍�*�W�:zT�JLjт��9�Œ��qڙZ2�q֙����|�ω{k����Z�e7���U-���]��A��AĽm��pU��Us4�����p�*Gг��o5P�i��7atq�|�R̳��f�Ɍ�c�D`d*4�w%�rE8P��ڬ�