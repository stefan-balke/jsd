BZh91AY&SY�R� �߀Px���������P�㐂ᡦ�	E)�SzS����i��1`!��b��M�OԀ4      ��j4I�y �4j4�S@ �A�ɓ&F�L�LRDCF@&S�M� 48I�BZ ��Id+��~*��C�]�R`2����m�t� �hY20�h�j�F�2H�������h�[8vC/ś+0a��2����ൽn���%�T!*���qȇ�1����}�r�BDX���NpP�-�oQ��S�b�y�q����`��n�X�}Ũ�Q_������ںL`���ǛW�`sm��e��KP�Ck�B"�Jl���V�Rh��-�-�Yf�.��ƬÙ�:�h]f"<��\�52��xj2GNv���ya
�C	�PTq��k�`$�'
e�5����Va��Z/���������%ŗ3���׃lZ2P��.�b�ݡ�"-![��8�($��c]{T�khw�eǘ�>���$!���m��Ax8�@��[x��B�<'��R�2��
��d�A�V�L�VB�mKD1�`D.� ʨСlh��aس���6����%?�se�Ѵ�nB� `|c��|�R�%���m����z&nk�7��U6{��^^>
�5X�s1R�@d���/��H}fލ���?�}��4v��,j8��r���;�R��q�-0�����>>��Cֆ��5ә��fgܨ��,��H�R���'��K,�3ߒV�K�z5������j�D`Ww4�k�.�K�T�FM.坥�w��N���YN�ֆ���dTn6.�S3-J�����l8��s���/��=��qJ)�����>Q�ח��ɹ�ζ��,1���z��YM������P��؝;*���@��E� (�)���ϖ^JUF�����.t=�/8��e�+�����v��3_p�CR�i]�ej�5�y�� �@ QåA �!!�P�Vb���#�"$�1!�$l)k��֜OFؕlx��s�ֳS�Ԓ�G����S��������=)��+��TM3�y���+�j�GYJ4�r��aX�<Sy��w����ۑ�b���)�κ�I�Z.�oÃm��S��w
eh�|ݾ�\�P��X�	Q�L�q8� �h6;3v,��.g�����ڋ̡Eך��/�R5|��S���K:�����6ɾ��m�c߻��|f9��i�P�QQ7�^1��ܑN$��� 