BZh91AY&SYO�� �߀Px���������P��D8���IFh�O	<�������h4	@��(�54  �@ "hP�F�CA�h  1 sbh0�2d��`�i���!�*H�$�S�<��44j=M� �M6��Er���3B2�,��⫵&�K�J&,Z��W2��?m�s� �4,S1a4wڪR1#'�a���j��/�np���㆜�,�i�N����c��Y9���n���Kf��SJ�������l)R�l\c���M�R�t1�ԛ5� +U�B$��_Un���� ��U��o7�����4��Wk���b2[�	��+[7/���r*�Ъp�\�~�®��~P�1�Lz9h���3Q��1b����F��������!uj/v�S%#������$[3�#���mB�LP��R�R�*R��}q�K�',�3b�U�[ͩ�1�ì����\�ߺ��e�!��f�)0��*9W��ͦ7��61���m��Ar���@㤶�ʅ w��J�Iv���'F��Pڼ���,F��{�GIzH�e�P2�B�QA@�5�C;,c �&���6���<�O���.�CY��q�W�8qTréU�a
{�#4G0O0K<�ǌ	�A�#\�Y��3o:�ZS����9 �lU�[������g�R�hX�izk����LҖ���t���I���'�Db��
�*W�6Ӄ��1��*W	��4Z����c��qJ��Ք���`�F8d(?榮�����7�X�/�U�9��1VS��d�:=K"������dc֮ᰯGs;{t̗1_��w�v�E!����/�.=�}�X,ߌTf�7ׯK4�5�C����|�M_}���!�F�bŵ����j^�m�A��2'T8NI*��A�ipTyX���ߘ��6�d�)1P���H�7ګ6�/m� iXX�ɺY2fP��\���G��H�d�7Fb�0-���bE���[�w9x#���r��[�
m|�Rd�dw�wg6|[^�����컛�+���|�t�%2�z^3%�+��uQ���L!������u��S����#Y��U�O5.�3U���f�5p������NA�do��"By���(d�u,�8�R��^�V���hӡs,�35�4^_K(\�^ُeHǾ��xjJ���������d�41F�ŜyX�r��h+P>,�N2#!G)tP��"�(H'�
g 