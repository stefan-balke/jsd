BZh91AY&SYq�rD _�Px���������`����h=;�:  P����Ѡ  �@   	M&&�$��OS��M0��S�4��	����F���i��&L%=BDM h4h  ��s F	�0M`�L$A2d�!2)��T�G�� 4(��ka+�!i c$�9	d+���j�bC�heQ.�"`"���_�
��|�H�U4�tY%G����k@��4ח�w�����v����+kH���6��E��.��8�`�	��逭Y!s�K�p�t�Ҳ�KM1���D\��2���B��$���7����F�ՠ�m�z�5Cd簱�&�pv�2]�����U�ڍ�}l�p����1���u��9];WV��c
������� �y�* �E��}�8+g�ZB�D�N�!�	�ܒ���|���!�Cp��p�~���89�ʆ���LC4�ؕ+��9b7��y�`d��J�ecLI��3`,H��M�*��=CJm�֜�6b�3!�D��ٞn�D�S�cjfDTB�KBy0���z}���.���[o�F��L�4�Cβ���a%1��<��H�\�ӬP�F����QS�PJu\cg��6:4�ˇY΄#�REP��d.UC
��rjӓToY�Z0���6ՒtT�ٷSD4�j0�ݨ�.�*�G+��8�&��ĕ�s�|�*�,�j�p�x�yE���;Bv���w{GO�;����IA��jh���ʊb�.�l��%`�
�fE�Q�L�T�fe1M���	B)stP�vX��*CM^�

%�i���@��9'e/��<z2�)�.�E�@@�p�Ǳ���fl��$Z�
� LQS�m���CE�/�Ć��!�f	@EE�e8�?'��t�)���B?q�×�����H���E�c���{�_Z`{�Zn?��k#���3�u_Bd�����q}11Jr��|��Z���$��g��e�z7$DU�Єpz����g
Z1_�U��Ċb�Γ�T%;сSU����"�xe�*�|�Y��?r�UJ�U�1;��y��:�姊ohn�%�W�����;�J(G}��b��(��e�4p�`���Te�18קLg#�`�L�5}���6}8���߫l�Q,[d��5�~Ye����SuDN9����8��2�+Ψ㉩�n�f�0�C����0����Xn���a$Me���7�"�+���Z�TG�[�K�]j䦅c�6j��{$E���[c���lJ��D�
m{��]H�_������K��ݎ�������7�%1�y9���ᴊ��S�ϰF�0~[��o'���M��*���:)u*I�Z.�j�_+sd��{S+FZ�z�ms���da/Zutb#&����ol�j��&l�yӡs<�G��0��a����v�r�)#��k��n�]D]��
ke�x��u��v���t����C���i��я�rE8P�q�rD