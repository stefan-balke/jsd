BZh91AY&SYR+ �߀Pxg���������`yî�� p)� BQ)�Sh (44���  h4LB�4��    ��L�i�����a�0  �IHM!�       2i�# `F&��4� �RDM2d4�d Md4 ��&�	!]�D�"LA3",�~��Xo݁����M @Lg�]��I!�	�M�P��a��l l�6�-���vz>�Oļ|[:ŋǋ1f-�Ǐ1f,�31�,ř;��xr��,7= 2���~UǸ�p� �;,��}���j�к�u�Z��Vֵ{UK�pނf�vR(�Bd1m�|c��*ۨrG"��)
]$���Ē�P9����i	�R&P��3>ȁ������ι�D�����Ҕ5���[�N��a�h�ff%���9�(
�
-��>'!PUS�����k�ܒ�	�Ht+Q �`���r%��F�y������Eu�b�B��낍�t�v��л� �M|���[�*�x�D���(m2�7���kLn!7p"s�	%h��� ��4�Z�d�b)�c�ȁk��3��yB����4$�Sl �ј��Bձ�R��za���'D.&�5�3Ll�ި��C�]�[�1�-���:��Q�͊��Bj�"bĆ��4���n��g�����q�r�n���01����1B� N]I��#da	�l�7�N��U�25��5��,LÜi�fh�92�����
jA����d��#�d�A��N��b<^�k8w���|֘�b�:�]�����S�3c�ی�Xz�$0��&݃<��=�Yj��bZO��V�O�u%���k����m�#UR�j��[��le���-sRt���B��y����d Q�ө����f���NX�(��UV	�_�sz���;��)�GU�ar�n����I��`[QJ�X�8�bW��-b�
�E*U�7Z"%Q%f����,h�"�E���%Cn��4ۆ���RAb�"��:Kʿ�]s����ݸ �>���p�#bV������>_ O0I>7{$*5�p��9�P34�i��L̶�l��{9	�phT��u��ȇ�����O����<��;�?�б�kx��C�_2bz
Z.=��M���S>�'�����N��Eݛ	R)jobz�Բ�k?4��b_,���2�
�Bs;��Ugif�Z1_�U���Jb�8ԝ�P��FMV�+K䥽T��*��盇m�
,UU �	���`�įP�+�OsCl`�1_������n�EBw7�<�VQ����h���fM��FXc	Z�ђЙ . 4�H���hK�}��V�����,Y-�|7���,���s�G$�I͗D!�񼢣��}^�~&�a����"d����e�0�q���ۅ���Hְ�w^�d\�]YglV��Z�>׍|�dk/�)�f�a�&Z�#K)���w$y�Į��C��H�{mz6ėQ>7�h>���)a��gC��-��7*%1�x�5�-���)Gg���]���m�]���v&8��
�Z�N��.�)I1�E�mRI���Y)ß�"ehˋYZ�68�vl&F��WSC&��X�rNCZ�����=:3�Bw��f��B�ɂ�u�s%H�񮍭u%"z�vv��hp��&�P�ot��㮪n��z?JmT7��)LOo�w$S�	e"��