BZh91AY&SYW�N| �߀Py���������Px�f2�0�S�4�&L@ �     q�&�a22bh�A�L $$ ����z�y��ښf�L h�I=&dɦ�L����0Fh� Q&�4h	�Dѓ
4�6�@ h��!>$� �Id�A����:�4*E�e5��͸m���в�4w��D��>n��ǻɻ�xwv��b��'N��u��-��;:cn�j��Φ����UzW��&�tς��2�6�;Zn�-5�C�:&��B�>[*q����&%���_��=�O8��S�7��xw�c"5S�����pb�T^�TZ�MvS�]*?�f0��l��h8�#��؝�ʀ��&|w)�k0<�ڊF�+T��c�f�a�މx�n36���2faH�
aOg箪�g�uZl��`��N��p��lc{m�����/�~���#�
y��*Q%��N^�i��LmbF䍍JH�e�4�eE�*�� �M�]�r������j��J�� n�\��(�����u�ٔ����P�ᆁ�����T��ZHCj��R2�(jIU ����6������i���=� ������6#�Zu��l���m�G�+�DG�k�/�Hj����R�K|���1Ilp�w�m2�I=˅c�}���x���E�D\�]g����|,J����Ur�<%�f�%��h����i�k�����I�˴���G�ar������uj�$s�mYK!��z:.�2m�*�m���ն�{v޶7"����1,<���4|�6�Ÿe�f(S��fN����$&#<h�C]�ǳ��&뺓�2l���4�f��U0h�-����5�[)z��AB�6���-X��RĄ�h�H�j+a����0Y��Թ
VRO��[����6��D�z���*JU����Ž�(:;��r�f��b|���%oC���dT�	�A)9�9�J����3#��e/GN����NK��JavE,�SL!�}8.Ko'���1�3s�J�-��Y9��Z.abTRO-m1�И��ֳa�a}�:�٦�`�]�v{"��c�=�[&"Q�(��mFi��F���Q�\8����3�-�/�-I�k��!�YYO��H�

�Iπ