BZh91AY&SYj�V� �߀Px���������P�:���	D�h�I��!����4� �5=	SOS`L 0�`	M5M4 @�  4 s F	�0M`�L$H FF��FS�6L�M��4��=&�'�P����$�@�>?��h�B
�)@L�5���p/���B�c@��jR!�	"Ȁ���:q�1�������|��7�@V��$G�߅����p���X�cS�l��Ј�G�`~=���a��@"����с#BzK𑴖D��n���9�1ZއlЄ����A!X��n��ac&�\��__�<�
 Ci����A���.W�,�}�B�(��&&��4���8D�^�6JU�w��b��1Y�	ZPq	VRT����UА�0Ff��%BȾ'�,\���jA,�dL[%�3�8�jJ�f�V��"�4Y+ V�(�!����UWSaV�Ś�8
���0��pB<A�P�>ږ�T���n.�b.̒D@A�3B�ĒI@��I6�����/����gm���u��$��K"TT
ZX2QH+WGA�H��22d��CA�[dIK��	Q�qP�BP[FBYut;,o�#���	�� Lx_l�>�)�8�bGQN,��n3�;�$�z"}�߽���w��8����0���ƨ�+�b��@93���+���?]�,D-�0G����~�^�0�B2�|�����jK˹�y#&l>T
	����i�2���{���i'�U��dTm��39�0,j��P�+�sT�%��Ćt��5|R��R=��p3Ǒa�]�@�m�����3�c��>����%1@P�a�,�Ht�3Mѐ��6�}��'z
�-	:�֤�zaUa3x3�7y�Gȷ=&�M����"4�-��z�Z�m�V- g]���ô�����l3�^r�Ցi=�X02&������r���� ���Z�	�:V&D4�y��T/	���G9�&�h�z��6A��mN�'�y�=H���ʈ�(��<̡�)I 8
��1����:3#�c�Ƅ��>��XI�����@�Ov�F�������yi�;e�p�%P��*6�3�y"��!���
��ѿ@����i7�"�u	�;��(�|���fhZ�A�P7P��I�G2��b�@�D���K��c�}�f�� ���.`l"�b��FRDw@xn���mT�e�dH���M���ܑN$��� 