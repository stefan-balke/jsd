BZh91AY&SY�ld G߀Py���������P>ws�88U $�5=Fi��i���m54d@���2djb��M       ��%=OP  �2� � ��2b10d�2 h�00	�G����jjfP$ �i驧��L� J�Aa
����[�|!Z��4�$א��m��4%�hVL���#j +l,Wt�uq�jc�o}�Yc±�1`!�)
%���<������ete�у��|�,�����b����Ċ�F��b���5��̌ M��ɴ��"Ց�l4$�S��1��X,\��?��j��e�P9$��Lwn�p�OC��H��D�4���rTP��'O��Cp�h:��]-{` 5�/9��6�XI-�H1
&� P("�Z�@(�I"�G7*� ��YR
V��#�:��kkV�+*	%�D�Yi�RT)G�g2���"�,nP��j����Z�!����� �Aa��J �m]*�Ɉߴi�$�S�#�#uJeb����J*t���)2�X��(I�cT&�����a��I	˅W7Ba�d��Y7�[�Y���hq�0�}�~��l��su��m���^Ro��b�+ɠ��&#��|�ӓA��C��b��-���=�,�5�}A�~��J�0�.�tgsWp���$H��dS������]�Β��i�6$��7�ʅD�`f���4C2(̂ޤ��@�kk��;����l�Pd�E���|qj�e �M4�"&a����v�gU��g�"�i�r�N�Wh���u\��qQ58`!�s����02KT)�GEQ��AvY��	����h[�wߙU�-T��&�c���}�7�a��Շ��pp�k�x`>jֽ�f�Fŵ�YW�K>�����`�-�T�A���QL(�0.(ZS��-��.&$� 	2�	�:V&D4��Q#QPa*���s*M�P�ʠ"l�Æ+��	�Nt�a���|� 0�m�{j1���a 4�ܼ�f\��k�o8n+�r:Ā/#��h�0f�Ni+3����8S���k
�4�BD&�)���%������XEp/X�ZE��&��_�Q%R�( g1�k�eJ�q ��.E%���U_�O��6�φ�{I�� ��d-Lcr��X�g���k�pT�߳1�V�����H�
xm��