BZh91AY&SY_��\ \_�Px����������`_�(5[��P$�i�'�mM=�     5OOQ=2)    h  ��M  �     SҀ�<���@��  �4 �&L��L �0L�0�D��h�L!O�B����@�4�S11 {��U�?��9gl�4)A4I���Q��IF�Q�a 4rjM�b+��n�	_6o��=Hh�˼#�G����"
�^E���zٮ;��I{�¯M�{�!ӻk�;7�̳��u���=��,�fI�#@��nRE��[t��Ia)�d�֜�\�<�s AaRRV'��e� ���Y'��.�3�c���]� ��<��T��=��՞~
���{�'giۥ�]I+
����QRi�O�tβ�V�j�a$��ԃ�l� t6C��B	z�2�5��b����ZN�ʪ��e2������2b��Ԝ�4fҭ��k]Q������6�6kUr�5�ɲ��\l�9NF�Ȧ�빛�lgW����aG�!�l⬑��[#D#F�M��L],)CM�k嫎���ʵ��/��S��͑�m@Ҍ)T�����MT,���#	����=l�b����EzUU�A�3A�B��C�A$�H���A�(I �@��R(H(Kh��o)<�f�!-
����@�"\j��ŀ���`�!�n�@�UB�q�P9��+0�& �9��� )���:<�񃋀�;%&Z����	l>nH���z-k���DD�N�J=�P�̝�MB���k��Q��Y:���!��?��u��*�d.'�k���yޑ:q^#6oIZ ]��3ƁD���ּ*�����f��`{;�x�*���[9�A�nUg���r�;8�-�Q!���ܚ�s�`ձK%[$���5��4tW��QU(�`P�5������`he��I�Ц(
�>����D�(�::(J2%�$�G�ϰ5�$A��h�)�k|�1�X�)����o���7̮�3��ܹ֦
�>u�����,�f(b�_HF����r��N#�9@j�e:�mA�q0��Nfd7;�� V��U
, �W
�Ɋ��Z��j��d�Wh�|���Idͳ ;6!=TҀ8���������P�\`�� ���'1���T��5	�t��! ���CE���:� �<�YJ����C�Yx�-�,C�p�H�dö%�!��c�`�y��+!Z�}dT��E7nnr��iAf9���P)5��`h�,�$��:����J��94�����ZM�A���2��<əVb��� ۮݷ;k�s*V�?�m4���B�p7���)�����