BZh91AY&SYD��� ߀Px���������P^�0【����=4F`�CF����S&�B�aA�`FM4��@Jz�L�S�i�=C�4  @�@���&L�20�&�db``$CM	����ji�&OS��4 Q�<�bh�	�*$�P ~?��9��b
B,!)�c�j��A���0���53 c2<;��޶�^o��{�8/'��ΝT�yw���rn��7fAr4ЊԜ�N����]c/�{xYў
�r�9�ay#�bF&S'��e��؃B��xL@+I �_���Am���Ա�?J�@��L|p�8���cX�VF�}�	˄�&JdIx�Gr�*�Ye�H
]x#���$;�H��agr뤦4r�4�3�P�t�@F�* iN�S`J�89���5q�'������5�MD^�,B��A�h�|��ov���#�@Nfa�"Т(��UX"I6��t<5Ɔ�.%h�����ʹ�AMZ��&	53���+���\a���I�4�q1bh���
%�ړc�iŬ�����d�s&�t���}uЬ��
�#h�Ҩ��g���n�P�T��<�FҨ�i����-�f��w��q�l3�9ٔ���̙�C�|T �0���{y��6�k*�� �H<W����<�[rD�~���y�^���q�LL��Y_�r�b�T=�cdx��Ģ)J�M]�5���7f���E	r�t���#s�0o0k�aIV8Z0̈��.��si���i8�_]氹���{p�Y��=2U��q>gxj>��u��H�%̒7�x]� ����(} 漂P�'�JP��cM�ar�t:G�K8%�q%� ���	�p�d�s�˻>Єb������{Opgic�a�@��K��)Rh*�'5��s�r�ɤ+�Ve�8iP"ABb�DAqH�\��}'q�N��"M��	D����{�P�E6��o(���]ؠ��p�'�F`�w:�A;'WH� �n�A�CBe����-�N�1MA�L��A@��d�,z����]ʡ�(6�E3��� �'��`��g�qa�6n�+B+�7`g7cF%���@F�,������%I;˃�Ҿ���r),aQ������1�z����z��#XL��c�F0��V���1��z�s�7\֪^��E�$\R�!���)�&�