BZh91AY&SY�F�� b߀Px���������P�` K�,�Q'��&$d h@  ��A�ɓ&F�L�LB!4��L@��h�h�   �A�ɓ&F�L�L)�dɩ�Hi�O�OS�z� 44�2yKʔ�U�ֈ؂HB?�?̉�A/� �B�1"ē)��_����H�ѱ �BB{!�L% [% ��z��������>^�\Kxxv�lg!��D��<_\ˢ/ЭA8�A��x���D���#/26���R��$& +F�'P�IDXF+E�/�b�L�L]P�ݠ���b?ȝ		�%������8�7�Y�F"*((�]Ӱ�	����]�����[�Ԫ��x-UŇ`m�����0��sV��hz��+0z��7��](6_T`�`��C-��3CDc�6�jp�� �LZW[)��fJ8�r a�7N�Sh���F7f�Q2`g���^L7��U�KF�S g�t��l�V���6c��&��0�\�������ڢ˾�F��ٌ�ն�gٝcG0s1���`�d�W���f�:���:����:`.�`���h�e������7��m�4��=�l�|�椻{�B�OߢT�K�		cÃ�(6�ۚ!1�668mjF䍌��# ʨ���PP0�x�3��ƨ�*�
�DJ����+��	�p���ã��>�Q���uF�x���cDԅU������H&���6�Վ��*�xP����Ț�z�Q%_�3������/�=��@��BA�^wǸ�5��5��A$1���J��;�������B���e#q�P`� ���lF	A��>�$H�,�X°�)e����;�/,�F�$���t�CZ�V	��
u�k���Y	�=����G���IA"+�#v����r \3\�����ng�����0+�0�M�&�(����vo*$=B8��r[��/
����I���xS�KnXzn��	����2�)�~�LaDיnb�\�h�e��w�������i�H(*Pb�{�Z���B��@����� �d��`a!������̎�2Z#FC�d ��W��'��F5��+�p� ���Rd	�?+���y���#i�< ��2;���`���p	��P+	� ���WPT�G��Aa�w����HVD1Rt� �)\I&D�F��̡���I)pgp��2ªL�E�
�h]6	A����zHw�n�L,��Es�Mh@d�����
c��6����&q�*�fXln(�i#~r~w�>f��-���ZId#-';k��ܑN$(�g@