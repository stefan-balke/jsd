BZh91AY&SYO��� �߀Px����������P����ɣ- P(�z4����Q�2= 4h 4���i�(        HHI6��0� h=@  b � �`�2��H�!15OѤ�yMM �i=FL�$'��@"�H� A�����I� �B��Ms��͸�CB��0�;��&�
�{����>1�F��W'��_6tz�Ơ��2d��p��;_mU�W$<�'&6�&�)	� ��=���}�̨�2�^A�{�2 ݼ�7_�9���h�x�BJ�;�0�Y}B�'��ۨz�"�>��#���q	0c�?\��;��Xմ-�[g�*v8"�.��T�;5�Wв2f6/�.���{8
�:��U����5hfi��F$���S�
`��0�L���vb"�(b�I���
P8��*]jC�T�8���A�� j.,�J�{�o��E�f&�w��R�*Z]PT�&�W��� �,ذH�\.y���fu^�0��E�g�j�Ak�{ѱ��o��m�4�rX���gx�T)!�rQ*Q%��:��F��k�ޣrF�<1Q,���x�b\l�ժ�b�
���� cCbϙ�M�}3ˣk�ܜ��,�;�E��0���Z�CK�'���%s��*4��Ya�rו��F{��sJ�1`1�f&�+r���:CU�kp�np�$�� �	�S�A�N�ں( �����C�x������ҪA���4'��Ǎ��3��!�I
���� �)ܒy�%Z�~���ވ��q��MC�ȉs�Mo5t�\7�o&��\5�_V	��C���83���kXw�!�4�
�B�_�~�3����q��\TS�=!���I��˕�ɯ1$`��Xlq��#1��T�7'�L
�L���aC�3���E�i��H�~+k �%����k\�oCK:B@y8	�9�G"� �W(��(Pȱ.�X)����]�Id ̀@����w�a�!/i(�E�HZ��2Pn�V�qSF�,�� #��z�M�GC���5�H�_4��b*�U��IVALl��g0�4&W��;ĒC�� ��Q��$hH��֯,t<���+��/�*6�3��d�3r;�ZD"���F��Tf�sa�3�GH�%"uPN/ð��S	D87��#P)5�P8Ե�$��:7I^e�Ր4g�T�i�����M�A����R$Xڰ*9"p� �xjmx�-k�vk���%����)�~G�