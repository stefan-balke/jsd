BZh91AY&SY��Y  _�Px����������P��M@�8 4 �MM?T�OQ��A� �  i���jd �d  )�������4�� ��0L@0	�h�h`ba"AL �$�A7�ji�22 =53SI4�y�%I@+�����"��sL���� �$�?AɅd9l3+X�h�ԤC"�"C��9g��ʎWv��cyh̬E��3���0_�O�	��2�<�e��*��"���n���T<�Q������|��a#�"�'����9���3-;� �lx���IYm�sBC�j_؍Ąą4�[��BeǗ%�h�y2�aui�<��Z�o2:U�~�5Rc^*�S�i�Ƌh��2D�?P�J;uY�fr��$��C��I�lhcL%�iFl��1FT��f0U#[.(��5%�6 �Ʃ`�0PIL�n�IfИ���Q�@f�T�Ё+,��&�M�wl��>%%��5����Vz�!�L3R�2��\!���(+CE�a	ť1{�u��m@ĶB�l��£�6d�]��L�!%��y���$D^r��1I'��!֢6p��I@8�*&����2��*����5�jL���0,e2�2�*�D�Gq,bP�I{TPP!,i���,$�w:�1��<$�Q֛Np��"Ͽ�A�{ d7�H�ka�(�K9���!�8i�޺ 1�'�'�����`���La�ڐ���u�t]=��}%�Ra�_��MDz�~�(* d �;�z@��k�f��^�TUЗh��F,��
$����%b!��C��dw�I<h�mѨ*�ka�X�j��EwK6�(%�\.B5tR��Q��g]t����e�GD�i2(r�o<�v� {�mE�Jb��*O���ꚧ�@1��(�!��đ��x����$A��h�)�n}6�(��
k�&r]����*Y�+͂��m�~%۰.U�pݵW�)	 ոB�y�@Jy�r��@�P�#��	��+��� E�#�JH(,��V4L��{�+0�C|��4�Ԡ��P�(ScS~B��B{5k���`3(G�gm����^��dM�q<�D��5�	��=aa$���r>��A0&vd��!hu��[xPm;�3<�Hc��Q���̠ͻ��U�W@gp�3�E��Rz.�PB�t�n/=�xԅ<y%�hq����,6�-H�E25b����L��F��A���|�A�	������3��ץ��u*Ye��=&�2H7��Ļ�rE8P���Y