BZh91AY&SYC�X� �߀Py���������P�]��0�+@	SD�O&��x)�jG�6��CMC��2b10d�2 h�00	LP�?Jd�a6��Gꁐ @2dɈ��	�����$H� �)������P =A���i�H! Q	Y����#*�i"b�����8" <��i*��GsLF-`�`�d��N��U�|��>�/L�
(x��yՎ%e�����:����?H��.n�"���d�H�;�e�%5%�De=�1Y��"�c2i$T>�y���)�����Lm�;h����GFu�̮��O/��kUę%~'F�������-f���!��H�5uB���)��s���ˑNy+�����������8����27P�e��of�XZ��9���THBBԒI*S��/�r�N�)]���w���oU4�2���WjHuG
 ���[9�YH�R�@��c��]�9�y�82�qt�A~_�M���X��Rc����9G�O@�7V��o�mO �܄���Y���е+8L�yr������/pB����G�i�b�(�� � <��V�+�2�R^��gx���:ͬ��V��j*T>��A�wZI�J���Ui:3��Z�S!%�|nj��	��DLj�L=��}	���26k>�*HT��~��^��@����a��Ψ(�b}�xx�tӥ0b�A���$�G����v�����,��Έ[v�� fS28�0���l|˵h�k2�l  #�2Ek^ͼ�hʳ4�Uv���;�9Kt����@�s���oUɆf��+��4�q���#�J�	�Wð���z�K�A,��
�0M�P�*M�7h�oBz�]G�̧4@0AF�Z�v>DJw �2�H�& F4&}<�A�,I+���a���*���>�����u�0��P�(6��3��D
X�"c�� c��ճvaV\����H�:�ԝ�o(*�Hd�+���I�Ɨ�y ���
K4* a�Z%�K��e2�onscI������0`lR,lXDw@�26��K]�38�j4+ى�u?�w$S�	>���