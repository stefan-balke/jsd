BZh91AY&SY2(�� _�Px����������P��\02�&����S�44iMI1�I�x� h����@!*z�#@  �h $$ADy4��ɑ�A�  4�@s F	�0M`�L$�L�d��M1M2Li���4�@&�IƽoI%�&B,�{����j@�0hT���)���Y����hX�b�$���:$1�3}�g^���|r���W��N��}6p�����0^>����J;DԒ�j��jچ�
��K:���g'N66��!���'+�a��jNc�&�|�(>eoF����(āЂ�C`��HXN��HRp�{}T����4�Vl���l��BL32a�����[�y�2X\-1��<P��ت�N�W'O��^4�	���.�6��Ի&�J���R�ABPy���e�Bd���r葵�"`�!Rf��")��0\�A
5	��!&p�WU�^�k�`��H2Ռ�a�]n+0l��`X�d[�	J�C�]�2�˰�$�J��X�+��a]���$D�2��t*�Mճb2�[SJ�;QJ0f_
�UW<���i˥�F+PN�m�ܸ�w�ٲ׌S�>.cX���7���hbJ����7!�Ry�D�D���ǌNU7T��?V�6�\s+T��X��$n��	m��.&Xj�:-�#[�t�L2HfJ�׎���U����J�j�s�DC�����/P�F%��dh��Ŧ�pߴ)P_#��&00�������*S�|ޱ�H�u����$�f��od��{�q|�?�б��y�����̘JZ��q�����L�I=	��'�5�7�	)��4��2�KS����R�2�I=
��Ӄm7�� �p��QCm���kj�tk`���2��0kb_�ƕ�6
�3����Ύቡg�4'6��9��+�5�ѣ��q6K����ۆ��Kuu`Δ�y�G���I���>�>1P�Bɺ2�Ei
.2+a��u3���7�2D�4j��,U����q�{��'$ׅ�7�������WX����9-�`�ȼ�H���U_��Ը��ab�d�(,A���{It��aX3p����4`#��d�6w4��q	��jI<�逦I,���l�W#9�,<�e�wD�Mm�{��9�����K�J��Ei,��ٶ$�_�&�O#��<i�׉�Q��V��(vնZ�z�Zѳ��ة����F:M�Sc~W2_�|��i��$Ŧ�,�6�5j�K�o`r��ђ�,�Vh�:�*U�J�;$c���d�2Fң�������9�(ג���;���Os�a�\_�;��C5����rE8P�2(��