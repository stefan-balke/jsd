BZh91AY&SY8�  �_�Pz����������`_�(0E�A@P$��T�Fh���ɣ�i�M4  h5O�@������� &A�0  �&L��L �0L�0�OHD�B ��    �&L��L �0L�0�D�M2�I��i �	�4� �D �����F"K�*Ф�H�BP��_�F����^4��HGkRrQJ�{���q���VR�Q��g�g�wê��o���������j���5� en�A��Lm�y�{ EA$��O( ��-Ih-S�5p4H!\���/����ޓ��c����q����F��15+��H��Db�z]f���̘$�<kzm"+e�F$�<����{���G�˱!&��m|流�;c��U�����7�v��ee\�X���2�(������<S��*zW�*���,(�&"R��JԉAu�՝ڬ��M�/`�����!,�p��"�B�ba̚K�D�2�� J�ŭ�U����2D�*���g4�YK*��K��c&���d[H��C�mq�$����`W�ֺL�Xۉ��MP�dY�RJ�r�A��x��@�yw��3��T��
�V�b��B�Ž����E�^�>�i|�0gdZ�Udag����;Q����i�α��l#W����Yax�UL��0��K�"H��'B"nB�dB�AL��+,Y�����q��N��H��04�7l ܜ�\퇏jk�Vk���jrqn���REB�C��"�J�)jYE�a�JƗYU��^�Nnf���\�@��6�$�����G0���s!Ġ��y�D����C`�Je4�ʙ_�L�W&��sT�Lp��be8d�xC�	�.Q(Xp��T�b[(
	�JA au,7�Ɓ&ҿ�R}�tf}l���c�S`�;�v�KqO��qc$3�Ip?{g|�Hc�4����(k̮�?W�{,�Q'b�6f[�(>�`�92�)I�%�KF%�Hjv�ƀ~�� pHL-Q�{S
 ���|-v@!���1=Ԕ"K*BZ�f���D��xT=|����OUU���X�������;5�B$J�^�qj��IX���2]"5|R��U��p3��X�s��@�clm���];�_ ���}�E�q���(y�S�e
��\��p2BT��* r�@��т�ka��"�QTB4Έ[�=�@jS^�gH3G���ȶ̴�R��� ���``<�j��z8�ޤ-K+@6Q!.�)�GQO��(�Ϡ1,G*I�����°��M�$!� @H��@��-1Ȉ!�?"(�@�%X �-r��J
MAd$�l`�2�ބ�g�!.Ð)��M(C�Hד��xg��DF� ����v�V���a����<� � I>�2I4``Σ�А�a@	�+���o/��_�Pm<3�D��8�L|L�Y�EFo�lEXEoZj9ZE��&��Ѹ�BU4Hd�ƓH`5�\ʇ+�\H.�`��Z�H��5�}�~V�������bY� ��!�	��PIq������8*Z�{.IA��m4)i.��ܑN$*@ @