BZh91AY&SY��%l �߀Py���������P��w�.p 8J!&�T͢���4��   h4 Ji���4�P  �   !)�M�=CM=F�=F� 4 �h�H�        ��!0���T���� 4��~��&C`���$�]��	�Bc���В�X��T�V �s���p_�@�%�̘A4��$i#)7��Lp�еe]e�]�ư���Ph��^Y�[VT�� ��{WCN��ɠ0����������5!�-�h���hp�-�Ni�r-�N�E�̭��剮m�U��D�h�z�I�`�̝IR��-��`y>��r 11���j/Fh��F��t��ҫV���N�^0��U��T�dϻ3R�ua�r��t}�� ����V�I��R��	WfhR�x�����$���l敆�b�AQkN�ZDM�{Q�/2"���d�r�Av̽�������,9QQ3��]��/1�=h]9���Ůj5�#EajÕ*Wf3��HBC�m��Mk��)#cQ
� �&�%B�0��tⴡA�W\�GR64dbSE�$�A��o5@��;+�b���u.J	� 3�Z�_�#��.���{%E�"8O	�h;��\�CѨRʢg��'�ۄy���Q���"L�$g��v��խcU,4�{b�Nz�c����=iǻ��u��g�;!��A���X�s<u�6����)hj�s�|����eL�`���d�I��m���0E8�8NۦRJ-N��<����
Ձv8�ͳfU�7<[f���,�KF���9(�S*;ҤJtȼ�B��1�����;��IVS��ɪgvZJ���fƶ.��1�Z��訮4��azX�s��O�݆͒���q�q�',c���Й���Ld�̕:DD��F�D� 9�R��:V!y^
J�g�7T,X�4|w�8�8N�&���mǀz�[ʊ���OQ����M�ڙ���#2���6Z`�ܙ��m�ξAq�H(-n��Ad�$$ �{�L"`gK��Ħ*���Q��2B�Ҋ��ڞg�$�~��t��ǣ�s��X,�����s�6%��䳗z#�kzoWY�RJc�y�%�V��%'�)I�������d���<��߇V	��U+D*r��S
�\�t9���g%7��Jb�c��К�r���%��ϣ� ű������5��-
`q��6eюJL.m���0�m{%�Z���]۪JG�Zt�ۓ=x��y��6.��<�{��U�f�S��ֺF�fm[���ܑN$.��[ 