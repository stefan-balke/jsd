BZh91AY&SYۿ�* ]߀Py���������P�@p���m&�L%M��	��!��h=A�!��@��@ 4   h   ���&�Q�)�Ph=&@h P�dɦ�L����0Fh� Id��&�&)��=@�  jh�XH+�$�Љ�"e����Uv�/dA��@ċ	(�����n�����Xa�&�;UD��@���::w�u�u��ñ���g���΍r�gL�xs~������Tm�~�ۿr1�*�1nI1T�r�{3���U���}Y]��3��
٣B���]����)Q����k|"8����H����HK ��<G��""a��i6�Ï��27z�2�p�Lm�>~__`z�.3mE�oE+����a"���R����#v��9���gS�+�c]�6�=,(d��ą�܋��p�mj���l����;38`.Z���Y݆����f�줬BF���5A-�
1biN�V�Y���uSx@`���Wu+t�2P��@V��&bS��=��f	B4Rְ��$)4t2rf���bj���D����I�&Ɔ�`����B�2[Uk2��r���n�q�W�u!�HS�u�=kE�w�c���m���!�{��C⤻��r�I'y�T�Ke�<R��F�N��:���@�DFd��Lpq�<fQ#��20���T#]�3�1$�9SL� _ޖ[xȮ�+�;B��L�s�W)K�䖭J���b�'�$�	��	�(ڣ���*���6*����ϥ�qD��$�p��y0��g:��m
"&�b�Jn�A򼟛1�R��q��-2N~��S.OL�I>D��9)��s���s��"���������2�±�����.C�����=�D\��g;WI2�St4(u�5��"������pgwa�Ĵ����eå�t�[@��R(HD�Aa��ᢉE$�{��)g2ӵxՌu�c�g۽��ڂ�G����*	���ZBk�O���슛���R� `0"~��y�m�+AP�&Yˌޒ|ާ�Tt��W��ۘ�z���lT�!���jlͅ��$hupPE�;�X����K�\�/�7)�����F's[
Q]M��=�+��jI��H�S[��Eԏ+��?SsIa��g;jjwt+��TJ{:��K�'�q�%EuQ��ܒda$��q2v=�s�8f4�*�q8.�L�-x�^+��$Ӿ�����Zch�IÎF��Ɇ&����X5���8���j �.��s,�$�f��®�l�����k����%Hw��u��T9��d�lCe���=�*�����)@��
�G1�����"�(Hm�� 