BZh91AY&SY�W� �߀Px���������P�rU# � �2�M=5L�&#��A��F#41`LM&L�LM2100	L�IO�A��z��@Pd  9�14L�2da0M4����$Hd�I�2dS�bjz�� �e='����@�IJ����9R�B
�)"`2M��M��čB��0b���JJ ɰ��3^��7�F��_\��ؔH���*�w�.v�k9BJ_Cc�3g2]m��]�"��,h1:�NSXE�2S��3ϰF����M$"��}( ���c�S��-^P B����>�#p���<�u��ؼVeVUu���P�ܾh���k�1/{.4��q�#N��X��-v]4�����#d	�d�X�z\�C����!���%6�AK�X�����0���kl(���K��I(��3b6�4�
��G.F�M�er��*$B2�YFM��HQhR��$E��$e�2�aѱX���9h\��w�߭ѝ$��������"��7�ֈ<k���ׂ���J��Z,}�l�$O�$��!V¿
"�4���fd�C���[��B������S�d �@|צ�"�nD����^�<ѓ6Jͬ���;!0�fT>��݉'�U�������[v�l�P�=����8&��JQ��J���*]g5l�<����8ȧ��^�����Yq���&P�Y���L�L��/Q$o�:>���v[���P�IM7ٟE��������1��}������[  #J��]k^��B��b�4#;n��� ��W�~��:�8k�X� T`j&�Nf��7<�(�M$a @H�֠D�c]�llj`� ��M����b堆��qQ6Da�#�rΜ@z���f'׊	G���N3H@��P�m;LN��5�	��:@�$����×���a3�%���z���Ws�4�Ӛp�2C�V$��0F����͛y1a�4����H���`�7~� ���A��bF���8WE�	�:JKT* a��O��c��bmi1|9� ���$X�^Ul&�w@|��h�6�Z���A�`Я���O�]��B@NQ^