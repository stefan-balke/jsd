BZh91AY&SY�T3� _�Px���������P�rlr1�
h:�*x&�4�#�h��d�h4�%!( �  M  )�"z��P��OP�4 4�0&&�	�&L�&	�����d��L�Pި ��� yD *�??O�r/K��hR)�2Mz��	�py��i*��J��em�Z�wu���Z-���_|�>[��L�5�谷�,!-�ۃ�+~�sA��ݵr(2����Ϝ��� ����^Wd(����.�bIV��
���2�&Pt|>m$�!���Z܉�
��z�~IR��ͳ]J�dg�;���1�U����]�G����eJn��$d����3A��"�"E�2
��*��ْ���wYF��p�Ȳ�XH$�M�Z��:(F�٦�A
�\���(Xm[x��B���IP���-����J�>�(W}�8���e��j�8�{eV��b�UaQ[P�4�2؄�yKC�d�aI��^ͯ��c��8�X�p��	�h���=ޱÉrSw��B�7��q�h	i�ӢS'/34�3��p�0����zx�Y���2.,��xw7!�1��\{���B�x�!�J�*(�~�E}%���2+H։غj�(&o`m^�i!�
>�A�f���@�kfj`7����\X���.Y�&��Q.�á�A�D���JMD����8���`��BC@�IC�`X��﷼��M*���.����M:S��A�����GÕ|��y �T4RSB��6m(���3�&t�6MUг����)H�ʡ��p:U���5�a����4^�0��H��x ���`����s�c�a-����hb��!Xnx�Q�1
� a5�(�a��;���ꋆUf�s*M�P�*�c�ߥi<rB{�bG��T��X���|����qx@<��\yd>��hL���fAa O���uv�H�&���*��1�u��P�T*O:tt�ƕ"C��]�2*3^ܯ������1�����BE�f%�p� �P2�e����KD@�V2���0�=�ZM.dy���H�س�2D���sk�ީfo٘���B��5?�w$S�	C:`