BZh91AY&SY��� ._�Py����������P>r٠0b��	$#MT��x�ȣ@�z��S��hi���q�&�a22bh�A�L %2A'��@�COQ�Cj4���L�i�����a�0  � BbCjhS�L��G�y � $=F$��! TH$�?/?�r2B�!Z��0L�^���n�1
�Y2�(8�L�7l1[:ƭz7��������+=ID��{�XԍV�V�$W��)BJVz6^�~��1��?�c��*2Č�7\/$`�a��fU`�V�b%{M� �c3ސ*�DE�R.t�Mߓ���d��p!%Y���j��:oj�P���uԘ��g-�G�-��5�+ص;�u�uJ}x��SH�ɇ�P7E
��v���3*�AXq8N�V��m
�KM��5V��V/�Ń5U�1:�ĵ�r��t��db�%d�5$�bUL�8o�а���9SpXf��i����$�J1�U+�RF��,�_�\�ܵ����0L�%IH?Ia�@���.��A�(���a����q��0L�K�c�ݼ�岾B����CW(Bї��o�}�)^;G�'<�=��LIVHS�d����*�-������;�9����Z�(��$q�i���ҳ@���&<.	�f�nǋ(���8XX<� �\&(f�.���ICZ`\��F1:�
�c;r�D�5�=*��A�w�$�J�����.S�˩�53!C�Ѫ	��ţB�\0k��MRg�&Λb�=�e�T��C$3�*;�B�Cm�jKa�P�z��*K�����)�>E �uuP��Mz�#�����ټ�&H�T4c)�m~��ʭ�Mx88[�'�#��1�)�'8*��2}u�o>Ԙ�Y�.]��Wa�GIO�~�(j�Xff\Kz*03&4�2�Xny��I	`0I�L2	
U�PR65�:��Uf��79�Ԡ��P�,%d@F���v�'�NP\M�fF>ሐ�?������ڲDþ�:�[�f��6	��>3�X��:@ֆ�@����
�AL�֯,q=E�����*�N�����k�x�(<��<hPf��f*�+xi��ii'P������a""C���1�I�
�EK���F����qtP0A@u����E�=�fI�� Ӊ�/h6�E���g$A��v�M�#�Rֻ�f���4,1.��ܑN$�=��