BZh91AY&SY�߂ t߀Px���������`>��>��F�__
�%Th4ѵ2�hѐ� 24 �jbi��        ђ4�h 4  �    ��AM�h416�@z��@4 i�)&�=������<������OQ�=@��d" ��h��6��d3P 45&jfUd�4�8IG���"���Y�H1"�I����ѷ�$b4+�.�;ڙC��γ��g4l���pN��������&�ހ�iID�u�x�sew�S�(卹צ�Ҹl��0�R%�0i��>;m%FXہ��3̃�i9�i��R[���F����A$�΅�\K�`0i|]�8Dc�G���;<J�`�i�7/��W�����dF{����\#
T2�rhCc"i�xغ�]�+O����&��2,�	"��ɦxlA=P�c	)��%�h*�(�Mb���T��y�"��j����3ce�ESeF4�$��*j�(�^��`u�qf{U�'-4"��ĵeБejC )CUd�N�h�u�@�Z�X�s%"�E%(聈$9���;PT0��0�iV$aJ̊�f0�k���87F�@�`�,���.���7�D^���1I��0l������!33�� Q@��SP�;"E���Q�!�II���Iq�!���;@/;VI��R ��HH!,qh�D�Qb!CD�)���g��]X8�Kz�A�>$$):����4p`L�Ep�#p��c������6�ұueZUH�&��f�1�H��% L���3h�����t�@\�
�BHH-F��dŐfB	!�-���jݝ��XU�]�"XPI�^�]��gʡQ3���|.�D�C8��� �/ޒz�k_�Xcc���n<�f�A����ٜt�T�*%���4�Ρ����P�uNhp3��.kX��Chb��WN�[�~ lϏi�9�MEb{�X~��t�0bK�Cy+��t�}v�܎⤭�CE���^R��=d�i�+�*��a�WF����3������Z�����K��= 4u�sa����v'����R��hn�i1��3P�m�����AC ���EC�3�ˎ�,Q�`�K FDg�jG��	�ȷ0��Υ AI��J��9`e�R��=./�2��ɑ�F�Q�0*ǌU��@W�(�0��)7�x��F��4�=v��i�::H�U�$q��|c�a��r�+B-�r�#Y��\���^9tV2�"�a�A��Pf�q.���"B�K���� a���>f���|vM�A��nX�R\޲,�Q?(w,�V=�l)�3i���-gv5��ܑN$2���