BZh91AY&SYRa�r 5_�Py���������P>�*��L� �E0jj{P��h<�CM  !�L�i�����a�0  ��h�C@=M�h   � q�&�a22bh�A�L $P#&��M�$�Th�� �'�Ɏ���BDD��H���}ߨ�l� �B��X)���f�%�,1������6��=���wofݞ��f�=&�|�4�'?�j�.��X��iT6�N���	����=��m݌J�q����L�ՖFCd�9On����h�����\JB@�&X_�n̤:w���L:�1�������-Μ;�L5B�H��S���[^�3���A�1w4#��Z��Q�[��JWJX���5��x�E�LH�ъZZ��S�}f���)jXu$�C(+J�;����h:aKN�F��TK�iVP�tǮʖX��W����@�w������7�m��С�`˴�K�a�P�S��R�2�$���H�$m�I���\t�y.A��F����1p��E�[��kc`�$S�a�]Y��8q���j�p�F]>�~#�h��0�_v�������Ʌ׏�$J@�+�Xhִ�_��gҰX�X�o>��0jfp�<#� �fg�6a�^��Ey�9��\u��+�ex��z�L�#6n=�
	����J�lhL;��a_:I�F����N�Y��j��&G�|8512|�ϐD����`�R��x�ԇ��Yc%8i	,k�
��@�߉�3.3S�y���?��`�y"��1r�:����H���8�G�M���ԙ#���.���8H���$���#�ɓU!(��a���4b�4
f�7����h�N��6L/:C-eO\Q��0�Ҕ��H7,�`dM!Bb�F��(,A�ybBB4�d�# �U����"#Eþ\JY��������a�$5�I?�>2�uJ8�N6˦ q��wPE �oAR(W�|�kGP0a��x+�#ᚸ��|���BCiށ�� �N�d�����q(3oGEH"���YƱ*J�%u����|H!#�`5Ä�]b!Z�]d��0��Թ���/�Q���� t�M�{AD����X�:7�={�m{��:�����s1=��.�p� ��"�