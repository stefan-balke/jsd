BZh91AY&SYfO�� m_�Px����������`z� �\
�P4SM	�d�M     O@
Rh4 h  �  0`��`ѐ��&��B!B'�z�i��@ h6�M�& �4d40	�10T�13T�I�4e4�&��M  ɦ&��J�","0D2I%��w��Uܨm z��*CZ@�Mz�E��7�RLhȕ�.��$�ZƊ��x:7z[���Ht�WUzΛ����Ļ����L9��OZ��D��~�^xr�|�@c�Kq���xo����tMuW
�X�/i`T�����}~ ����̌�GP�3��8'ā�}%�+`�a:��>$�K��X���l]�%��?�>�H�)�ww��ǻ�5Z�L|~~�F;�^��BDJδ D`W46LI��O&$ �	M��{	⋪��2aK���#��G�]��iIj����z�gs�䴎W�k8;'+�Ƴ��GO5Ȼ636�2�]D��O����3[)OفL�Xk���Z�x���J�7MfM>So�&4ƬO�.�oyE�g�m������H��c2X�(����pK�جN�&h��k*��ò6&��c�Hb%��U2�-
���+�� ���7.��ΞLr�U�����6����e���jN^�J08e ��0o��� kip�)��&�S*�ah�kC3ö`s�<�Љqyۗ��%]���+�ہw(UfJr����˩�rl��hk-��&����D$N�-���
�Y�����#�V����fʹf
t�y����26���o-8ߧ���5Z��4�-�TS 8BB)�j�Q�{���a�AB��PP0�x8���&�I���L�M��\�m��L��8@\ٜE�����X���W~k���c��n!˨8�w���I�����~I;�6ʢ��WtHη���O��K��y\ͤOa�����/����y���T���B�f��bއۿ^���R���^?����u<��)�ޒc&�e�!>1����	)�Ct��/��Z���bz�ie��'�I[0.�3LTU)�Pmx��UeR�Դ[^����
`�Ƒ�(������El���o:C�=^#G5���*"��*�Ql�G�i���^���7�#9zX�wc�;|3�9b�'ONԥ�ƺ8�^,}&���vQ���n�.�'\�w/q)��q��e͟+l���9�
U��]3崦���u����^��Bw^�;G=j���6�,�.�[%��K�ZB�٘ڪ���*�1ab��pY�X萌A�H�n0��3W�/ł]Q��e-}(����%m�sHN�[�0��%�#������o�͑p��l�ލn��*�6�%<�'k��q�#8*4�����Bf_�sC'��\��<X��������1�%���4��{t0Sw�T�э4I�ѕ�W�_.�x��,�(��g#�q���R��f��V��Y*��.�b�^���ʑ��Z�3o�*C�g������7�,P�t�w���w�UOs��,�?Zf�mQQ4�?�w$S�	d�\ 