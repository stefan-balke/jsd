BZh91AY&SYOh�� �_�Px����������P��8 �d�F�$��)��'��4 �  ��!) �`0� ���Q�l�MM�S@ ���0L@0	�h�h`b`�$�I�M6���i�ɣP4�� 5=M���$��D��"�&1!^���W5��DhT0L���͸/U�F�B�fXA4yڪ$bFd��u�����%v�{���9=��ٮ���pi��Q=^?����p�߱ݝ1��ttV�}�Z^�o5���׀���S1ǅ��@������8�0�1�9]=5��I��W���F�����JJxY�t����_�wݐ��2�!0�Ɇ����m[V��.�W}��	gDQ�E�/�����K�7i(M9��:Z<�&���n�D�a�jɘO��Qv����"�KA��;2@����"/x�HT%�[�̢�C1/����KJ:Y�L�(�p���B%A�J��=� �Y��Ih��:A��@�/aP��ma����r���,.�U�T�E�oƽd�C{I��4�]���H` ��捑�n��<��!���o�m���!���t.�9�Ry�T�Kg���H�a��]K�6IaFk%(��	 K�FFJ��=�A�T(P�h��a�[|Q	��6����S�~��َ�fxk��g���>���ą�~W-�t3��\>nR�'�����VR�n��>���]j<��w�N�L;t'+t��84��}����b2�R'�Z6�U���׹/7��,=��3��=.nN�����D�F�ox^_%9�sN���E�����v��=�RJ�yve���YT7:�Z�ԇ���Z�j�t�i�v1(Wh�k/��`�;<�ڇxy��֞���9Ƚ��baد`�V�9�Y0rK��ޗ�p��.��!b��r�$F	���^0�P��V�2'��U��wǫ�Jr�fa'���m:�f��N��"�X��j�[p��M�I�6_i!��D�z݂��̮�����/����]```o,��X��ۅ�� F��TAb��萌G�K�\4
Ã�3���.*h�|fA)fHoWwu$���t�&�N6��T��o����k�/m����v&�?���]&j�L|�S�b�D���Tj)Gѽi�<�KK�l�l��i�06��3�2��\�",;��8��fFt��X�ơ�Qm9f���YS�^��h�$:M���5Mu�X6i��i�A���"((9L������z%��(����Y�S������,�ˎ���{�/�,�jmT3QQ8����ܑN$�)�@