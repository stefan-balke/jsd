BZh91AY&SYG�� �߀Py����������`�j�ٻ�����<%S@)�mOP�F�@�=M�h�ShL%d�  �  2i�# `F&��4� �BD@��� ���  @��L�i�����a�0  �$�Ba����i�&���� �Q��j, Oh�$ � 1( ||���B?q
� �Mr��6�쐖q�b��&��EM�#;��r׿���7c=�e���w�msv�r�iv�wmh��5YVQ?;�W�X,�>t6;:cn��ؓ]��`�80ť�T�|� ��߀���AZ�Q���S��D��ȂddJi��Uv �lw��R�n�ą@�-A�bi�.��ZUS����U,Y�$Ă ����D�]�-P�V�'��D���2ʖߎt�bA��r�"�8��Qc�[3a�4�lM�Q��j��x�6۠�̥��0���Ħ���Ze�ޥs$�� V�Q�$����6^M�&-���(��e |%	��ӽR���X8҃���&V�N% �RV(�l�TG����$%S4]�GB�C ��+,���E��˘A!d�(��Yw��9���jat���h�:��8�{$�4a8��K��A9�23:��QV��S1������VŰ�H�Z��b ȆmZ�#e�E`�pK�u����m��T$���>�����7�m��đn���h^.9P��u�b:����`�9����5f�`���J%�(��L�Z�Q �!BS�2���-�*
����Ě��"*�"�&����c��8��z�Ѐ3�P�燥�հ1X������u�CD��B{�|�H�~���Ѷ!�gp-�Q���`�>��q�ֺ�����E�F��xB��/:�#�w�b�s!�^X �O:���1g�!V�{P��F�\´�����(T�C!��<kw��A�O�$�J��*ƇcA��l5j��DΫ����d���8& .��/�U���6���!����9�iܑ�6�m!Ʋk�a@��?�A�n��Xd�(+�xÿ�}�ؠ4$e�΃e�R:��g6������3@�TT�E����P�&B\����l��j,Զ1�/�p�Mt�1ݢ�X�%�r;��@4q'�?C�sO0`P�p&00*؊�2
ằ�Q5�� �F݊�X��k��{IE�.�f����.*h�<)$EL`�kf�'�ͨH���`^%H��;hl��8���ܺř���c��Be:E�BBH|@�E��ON�H�*AQ㒴��|��/<���ci܁��� �TK\B&<Pe�Ɍӛ~"�]�����I$)*�U;n�M	�Hd������/+�V�a ����nr��h�ڧ�i�=ؚ4�G��������C5qX�d�ͶA�����7)Җ~�2��u��ܑN$����