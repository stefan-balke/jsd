BZh91AY&SYjˮ� ?߀Px���������`<�n�Y%�� 
 �{SLF�M4 4�� d  50&*H�       ���a2dɑ��4�# C �������=@4� Ѡ� 9�14L�2da0M4����$HCF��I��(b`�@�&�����Q �$@�y�㭤6�\���
�ЌQ���m���B0�Ƌ@@�.���HV���'ܘ����&Q�F����&c��KD��lj?L�s+C���w*�5����1X�X����b�����	1qd`#Uc`u�r3�Z�U�fgÛ�FŹ�t�p�rh�M�@���D�z�$�"H�m�56c��[0(`�L����G���,E�~y�M´f�+
�9R�~+Jͫ�\�[� ���r:�Q�V��;Z=(�ɧw���!1�<up�a&�KP��a�^��^�"��	cp����<�[�ĕ0�*B� ��^����R��d�4�"���^m��2d���\�dH��c dK"E�L�v�בH���R��$C�1��BXRH���Fa����Z��A�@����j��]��*:�!�҈�%���9�61���m���6pw���]%�k �B��'�^k,�f*��Y�nʪlaJ��L�$�P�BF�	�H�HCX�-��&�M|cT���D*F ���ɂ� �F����( Aje�:��B��,	/ �$jc�G��f� 9�����DDDQ��k��"���VD%��#^�ų��? ��0K��0���G��-0�!w��@�@>�J�E��BK�$�K��"��P��Ł�|��4C4(�3 ��[�$�dT'k_��%�۴�Y�7�B]xǉ�td$sLK�IA�"`��e[B��s<u��u�5��X���31*���o�p�o�ͪ��P�>����v����y��9��U���!U�д}�q(��3�L��篧�j�K�Y��RѤ� #%�b<�Z�q���K[@���	zzϨ�����(�N�ۙrSH���L5���m
�s�x���	�@ Q��AA�2�	�^�$Q"��Nl�2ÜʓD4T<�D�M��}|���w_��9���yv$���6^FÉ x��p9#�F��!�hХF�m���:�������� a���	f������`1vv��i䁜����L�H�&>$�jB��:��ˣX���ՊTy�cqK�9s(	TȒp5-A�� �P=G:���H/q�v���(���ld���6|��� �u��R,oX�Ig��$r�@|i�k�rT����h44,5���.�p� ՗]�