BZh91AY&SYP ! N_�Py���������PXo1e���@� j��SF�ɠ0�2 � �F�%L@L�h�@    4 HH�z���M�SM   @2d�b`ɂd ф``(F�OF� j�����zC@2i�����d��I" J�A������A�B��XI���K6��	d4�1CGrT$`�$��_cG?O]��M�q�^��T�'/G�u���%OL��P�-���$�����e_�E��RD�Q!�����-s��r���2�J�P�K���! T��H��� �ah�2�(���&�1ݏ��<���������2�Z�U#�J��k���b5�sp2����M����y�����e�Ŭ�Roc��.Z֑I{���h�Xh�ö�.�[Vʶ�
]mT�P��Y+��) �V��c'0�'Ux��	'Lj2"�%�tҨ�Ĥ���+�Ki�7�lcw��m%�}����ʅ$�8�(�����͍՛j`;�Q�6�)��j����$p��#��[
((F���Ahl[��:o��#e����i��)��ῬfI�@A�Q[w��y$@��udsU3�~��HC&���Bc����_c�[Y�q�&H�K���>�����pq��AHfq>���|_"��R*�o%�ڼ�WrKϸ(��%�Y��f6�6��P�dP=���W�I�0�)[5*1���:�o��ȋ��vu�L���֚@����+*���9�T8��,/V��N7�
v�@�XbX`�qD&P����x�1.x��+��7�:i�0�$@ʈh�d���d���H�	��z_Ͱ4�,��bV�Y0 h^y��f{ѥ^��%s��8���S���s@c�R:��`h,��j#v�j�!,�
85("���$$#�K�\2
��3 Ts�RH�EC��$�<�ڄ�ǐKA�܉�ȝׂ��}Ǥ�,mƣ2����a���d4&wt�R)+�s�&��c�3�I)x+J����醐��w f��"1�K�� _���ٷv�M��`n�J�"�@�����ĨDd3J�F��i0�7ж�H��/��q0Q(��/B�kH����li4$�� ���(�5����H�����Ck�f�[>��A��B������H�

  