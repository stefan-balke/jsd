BZh91AY&SY�4�� s_�Px����������P~wY�t��
S@4%&�ڞ����<�!�&�z�4� i� �S�H� �@     	LR54)�=F@zi4 z� h��& �4d40	�10� I�$�S�*{D�<���(  mOD�I��BI*$��
����,�_AV�!��
	5��yLIh���TwD�]��rl6���۫�l��,�f��Vl�(��_�����b ~��n���ח\��bO��jޗ\�#6�\E̎Yqi�C�~���yDjݨ�)�A���w�!
�a}(�+���ѵ3��/����{o;� �F��;���Bd�Q"�ڐ� �Dh���QQk�b:�
�MJՂ^��V��x��2���tʰ�(�g��YY����0���`�����#­K	��0fS3:�C�2�*�h*DR���``Z��Mi�%pWċ	�*��B�P�!µ�b�"���Nnfn��F{����e�4��97Q!	K��I* �wlu�a��n�q���A���DA*��F!F��_�K��D\lE�҃Qʆ*��R�[4 @@�m��!QI�~����6;������b8r���'��S�QI��m�3wDy��Ѡ-�Z�|��!dcIx��AִnJSH�����Ƙ�����0P*�s�5��)��d.���j����.�%�*�� �G#6������M12�eñ�A�[�$�J��슴�`k:/���c!C��pj�2����4���!�W�+
J�{��](p3��X�h� &0�	�B�;����YH�	N��'�w���Sd�(�d(D�.���l��^�odʡ�������QnT׸���������>�("zj,@PP[I��d�d�z1Y0K1�`���%z��9@m�^iY�.����d�Nf��7>I�2'UU�`0��t�8K7v��D��Bup?�ds*M�P�* �� #��pB{�J� �6"�3#�$+�%	������o1��Ɠ�1􆡡3���6�� (���`�=��5 ��h,tE��Ws�0
�4��� ɢ�$Lqxw�eFlݞ�V[�<M(fv�bu	�=�(R�B�`�#P�y@΄h��Z�����D2~*}�#W�sI�Pfnn�3 �=&�q�)MJ�N��7�Z�՚��`��h�뺟���)����