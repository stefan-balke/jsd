BZh91AY&SY�s�� �߀Px���������`��� � 5L�O#Q�P F�M   hIM OP   ��	���dɓ#	�i�F& �)���h�F�     sbh0�2d��`�i���!�H�I�h S�&�z��ɣ�MO)y4	=�B!!�B��JB����F(�*Ф�0Bd���g��B�e�! ��Ԝ�!$��_?8����^�.�Z�S�����ꩨ�-Bֽ�TF�Ll�k�z������<&S' �K ���e��L�WYY��VElZH$�Y��>���=�auJ�i�sz0���wh/4L�(O<�Db�;�f��7[)�%P�%�0�f	/��'�|Dm�����������p!1������p��Z�qh����4�YJ�k&�.��dʵl�N���5��;ګ�a#� �"`K�q�j�N*��9����+��3WȄ�V���A��Qj��O"����A$�����AtB�F.@��p�	��^2��% �AS;��HgV����dY � vT�lB$5<��H��a�pK"�e���C$EE��X���K�(��i
E
�1AuBZ�+�c�@�&ޙt)��"`J�&�YA�b�#hdgFF8"B`��N�ΗJ
�W5/�T04�R��@��F8�e ��ʘ.Vm�C�844�E���X(]7cm���Mj".J�iv71V2��`�DAU+Ƚ�vM)��qޜ>���G<QuUZ(�C��9�!޺�.�d,�u;�K�I�i&�EZp�����wt�$�M$H�Il&�y��f� �Z�Ռ"�BB��L.��T3n�#\&��J�ZZ�Z(FV��9aJ1��nݘ��B������l*2���Ҡ$�K�;�;H <��z##U�):0��%|���.��=0(LR�$���/�8��v���?��� ͐���8^u��M�E0�B�br�^��5s/��7$��I*�Gx!y�&k<�6�5�+��P=��A�gRI�@�kf�܄X�M�GF���5�B\���� e�I���"`��JI��3�W���b�oX
M&�8ȡŨ,
��p{m�-c%1@P���;����F���/,�a5�G��篰3l�L�eP�IMc�׸�����g2�Lu��E�r��\V�4�9W���z+Z�nچ�Vv�U�]����B�#�l5P.9��o@P`bL0i�d��|�/�j�p�@��ʨQa�l`�!A�"
$P.	՛FTs�Rh�������s ��0�$��j�M ��pIL`}�����i�O3�p{�7" ú��֒���1���2��I�B�:��9:�A1@ߡ\f9Β��,��p
��� ��D*�	"c����Pf���a�7ܒ�o�E��Rv���!T�C �k0X�P�q�T8T��Il�tR��������M#/G��kI�=�9�AkA�A"�Z��A�H������K3|� �h5�;3S�rE8P��s��