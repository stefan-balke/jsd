BZh91AY&SY�-�$ b߀Px���������`?y�M@!˅�`��=5SL� =A�   	M	�J$jb`���c�A�ɓ&F�L�LBD��G��~��!�M@F����a2dɑ��4�# C �@HɊz4��?T�)�?T���S�@4zL�R�I �I%SBP"����7�.���I�P!M~��ݷ��$b4�4$4lj�`�/^gs�N���;���i^\�ΟH������bc����r�m�m������c���)�7 ��[���'��ݺ%FT�`9<rr0�LY9%��_��}�0Y;ܤ$���j�i	X4[Z=ɍ5�~�vՔ�BM��ӑp�$��Lyc�5���#�"�\��m�Qs�n�Y��!: �o�:*��+�t����S,����s<)V��[VkM��̓�#9q�
����+#�(���ǈ��!'/�+��`��V�#	�R-�
���m�Ӣ�nMa�E��i�X��s���]�}�fC)ks�k�Am�F'�\	��H�pU����%�F��D���І��'m$�3��;ƌ�8M�	�RF�Lq��&����S���U
R�\�+G��D�$!.D�I0�J�q~�x�.M�r�I'y�T�K]�/��:腙�^+��[�Z!����ma#d���4.6P�*4�aE����6�Z���}��IsLe�Աr ��?������'-�1�(:<:p$<u��(8d�}V�u�/�����V�gs��0��5B �V"Iz�}g�ضz�����:�$��Bӝ�;̮��h2�Y3�^������e�$�.�K�Iz#n>3	������I4�6��yw22��Od�4��N�Nƒ�:�-*�7Yr��7ںI�o�4��`m�"�MCcC���:a8��̜�}�gC��B�����մ1,0Rd~��=����0bK�$@�Eu�G
���;�ͺa2&ꡢ���ۻy5�/R-$pk�ٴ-�����!%�U�& �C����R�7憍������Ix��v��ħ�>��)��i�"P��)�I�R0
A�_(�a$$k (��PE�;�a�!��H�XQ)1�D��	@�������	�>�%�v&/;�Db=c�P��؈�Ǿ&e�M:G��	��)�p
�I'�Ě5�q�s�IbIL��k*XvXuP5\Nh��D�5 )ܑ1�%�8hLf[��T�)�4֑y�bT�J/V��bJ���@6�+�Ѩ �L4�]V
�i.D�
A ���ͤ_����h���SA�%��3Y@��@<����7����C��㝓��ܑN$)KrI 