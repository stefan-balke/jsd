BZh91AY&SY9i�� �_�Px����������P�0�3 �-j�$�ʞ&�hO !��4bh ��	M����i�&� ��hbh0`��`ѐ��&��0`��`ѐ��&��D��4ԟ�i=C��4�i4� Bz&�1	�$(A@H� ����c��m��hRCIX�2M|�����Ā�4*��a	��Rm���Y����{8ve.�>��;,�����b��jn�vY���
�)�0!MpU��{fů+�ws����=��RXE��<�m�4�F�:NL��Oi�D��,�l�Xa��ᚦk�m�u�?��	��o7�S�qɞE�d��M7TX�36t��
��r���Br�yj����G�\m�.��o9�&I�:$D�)�c$���3u��C�+{���E�tn���^`gL��<�}ܱ��aA{�n&�&�b��(�Ε��A���yE���$����
�q:M�d�!��:�>Z�L�=�`�{J���w"����7�2��_0ì��u#����3���m������L���Bxr T���'�$�J�,I��C�XP�AH��D	�^�@����yP�i!�0�M�� :n�eΘ�əmqA�߽h�<ĲQ6;G�xx׋�ʱ�b:y��}7,L{�%5�Oh!E�W�jV66fɑ�;,�Dg��g�.,�}���xZt��r��|�x���@`�3���u�a�T�"��7"@?���'ؾc7�Ҧ��B<�1>s	�̘�ƨV"��P=ކAyo�$�J��D���XO&�Mը72<ze�S�Ę,ؔ���1;��YU�뮴8��*^�sA	6�C�	��B�NC��{tv��i�����%������`�Ä��a�|r0H��1�]3������*���n���q� b�[	��)�9R~��A4ܾ����JR���1\���!�s�Ga]���8s�d�'xX���HpL%�Δ� ��p ���1#��"��t���L�B,���%2�b��Ń�U$E���e�v��Oj��X.5�D2G�\���*tD,\T\FEAzW��-��u��aRBC��4�5�u���
O��d��w��	���eL�1�������¿�3(3��Tv-���lu^�`���x�a��q�t��Q�!HV5�@骷MIj08�9_|�����NM"����{I�� �x�����	1��J �H������y��ko�̓A�b@2+���ܑN$Zi(@