BZh91AY&SY�pvb _�Py����������`�;{� � �SԚ�M4��S�`!�b�1G�4dɦ�L����0Fh� 	L�Q4ځ��     	M%OSh&�Ѧ�CM h4���2dɦ�L����0Fh� 	0
f�����2G����i<�䐐� �Hi$��(w��L#�hQCHR�_@�dۀwHH�
���͠d�Ģd��m��б$u�Q�+M����TĎ�h�W
Bܐ��B�N�8"�Z��.\}���0a�BI�NxN�s�>����{yC�mbLedd9��@�<�#��Ȥ�[�)z�b���$���JH �P�#�K6CF��[���R���8ʉþK���)����s���1�������S�;5�<^��WHʎա�e��D�8(S,�QBը��\Y�SQ�<g	�F����AFtʈ��3�֓51���:���A�j���vG:���7z��[�rj��c�F�(����}9�nr�S�yW�ǂ��r��M�$e��t���rЪ�C�NOۜ7QUy4�@M�Nkj�\X��n���#!�^�%c�f��Q�7
5�]�.��S�%�qѨ匷:ܝid˖T���ڀj)��TL����֌q�*[9���֌�����3��:��ӫ	ه_]�3Ta6z���x�$!*i$�a00�DE [����@ V������B1��Bm�� Bф��:%�L�B&��	 �ꨡE�LD2�!! ����^� $�!�:r��3>���E|��`ݗیTe�<yRӎ@0����p�����CH��g_����;8�.��X���&d�����C�;0�>g�n�1���Z\���f�A��� ��\t��߲�b���dP@��-8.�oIP�I4U����͚�	����*�L�6�[ @�5zRO�iMVMf�٪ ���?��j�Ab4!tx50C&%�4�dyD0j�N�Q�C��j\��NR�
Ρ��0��
t�� �Y�35����B^��=�,���ni�1�^r(ʨ�y)�����CE���M����I{I��|p�.��ו����ֶ�@�/�p�)��ł�pB���u ��O�~�����0*C�1�� ������nx��E$+A��Oz�W���A�;�,8��1*��,�P`{�� t���ےKյ	봧��S�/@�4�a��
���b��\��u$�������hL�)�8H�E�9 �@�˂��"� D���O)�jaj�@���s@���DcK�V��&?�(F\p�Tf��d*A�8Z���X�%@����B`"��̼�.��izV��rX_iը`�v���YIU�;�zZF^/vF�&� o�ƃ@DJ�+J!L���{ 
\ڡ�mTժddA��B���]��BC��و