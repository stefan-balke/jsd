BZh91AY&SY�� �_�Px����������`_�	�e���Ud��$5=OiMSCM�2  A(	�$��h     ��=ꡠ�   h  i�z�C�� z�@ �  ��0L@0	�h�h`baD�O@���	��z����  z!�5�QgZ�R�"�o3[O_�K ��!���ah���J�1�!�
Jb4���Xj�Km-�ݷgOf�pf��mY:=�ZӢ�F��])�u��t�\��Sn�����e7���eZ�,�D���;vaڭ^t�;B�ܵ��Ok��:w\�̎r_�1F��m���eJ>��K�Іמl��"fz�p�tc_0����M1���j߿�ͻ�:������~'ɇ�Q�N�_gxz�)4w�4��^�E�cB�ܑ,����T�i�aN\���N?�d��,�K6�u�vZ�D"M�C��T	RR����e,g"J!L����`//
%F\����CQ.*�M�Bj�������^.<��`����r)EF�� f�h�KL,���)�Ⱥж-���%0N5c]��##BP�̢�S�R6�x�>���Q�4f�9WKWUW�QcZ�6+��R!�f�H��ёs��f��!��J`�V"&t�Ć-f&v�R���e��T�-�!�B�Pa!J��.��&�QF��gF0����$�-���ot�8#��g6q�eL5KH�ح�74���{Vg2�Y�Qo�r����ΆZZÍU\��
܁�` D��zny� ��>�J�Q�W�b�V)�,	�D�ċp0Nf	&�*M]HM��!�<�Q*�*�� �U$T�`ˈ�n*>㯍�(�:�s]����ի��i��4~L��#b����l�.aÊh�]�n��3딄$�;o*����V��i�!�
"�X�Z��N�ϱ��$���R)#n�q�!s���Ʊ��g���c		�A�pTf�C�K����9O�h�!W�}�Z�O��/������2�E@8��9�
� ��0��?:�nAlc=[�aE���Aߧ93�!IY�[�9(�%N��c[�$�Yb�`;Kz���%�`���yĢFI$ �+y�vp���L�[�Ed�%��"xZ���+�)�ۇIg�,�p�����W��A�	+][$dXR)�)1|�D/�)�'���V�<`-l|���s��9t�M��1�Q�{�H;Lw�ߖ��hw�Ƣ�@8 �����T�o��it@���daY�@�3���Q$2��!�/sҢ`>3 -^AZ�w�|<��6.�	�$L8  <a�e�3Tj���E�o�*1<l!td),�6�`�YQ� ܣ�u�v��
=���.�C3���A�up�l�QY!��!1),K��,�l�]fd8���RcXu�)����e�m9��2pib�*�8���!��u��j,�E�+m�$ o�[{�&��hmJ�2L�\Í��!��V�����`}��]T=Z�}g',�~��D8

�gqٹ���"�(H|��� 