BZh91AY&SY��s� 7_�Px���������P>�lԌ`(ր�(���S�M1j�A�����&L�20�&�db``e&#@�2=�4  �d sbh0�2d��`�i���!�H� I�=	�2���SjzOP �hOI�4���H�"���FB>0�
��`L�������a1��� h�j��� �@�����;۸wq�e�2	�U3"sor�kz��o1[i�t�:�����oo@|6�t��#!Α��&�#q��-���>�,�.s@
ֳX4W��v8~MN�X�����>{�����%���s�[>��s.��K\�׺�E:U�d�/�SPc�Dk����=�#Pm4�{w�U����DTi���;�&�DZh�4�u���`�K7EcP��2�6L�x�QaT�Lڭ���ĩ[�"��R� �L��,�0�cV1K���9��61�m���q����R\��9P�;���XɬG#�62��P�{�T��"��.ȑ��20��gE�ŵ�Ɠbӝej��k2ǹ��(I�ч(84�f���6��	�g�$e�>�q0A�,U���"Q�ɓ�Y�V5�Z�Rhf��4`#E�.�}/��h��P1a�鸎�LyE0�B
��|��+�2��/?PTG��3f��2������d���Ԡ}]̂qoRI�J��܊����q�A٨5d"����PL��5И:DL�	R��S�.����!���5�li9L
���p[1��`|�������>��?/m4�0`��.�H�8�����&A�PT� �.*��� ��)&٫�%�GD�A_�ե�=C�Z׻~�4d�4���x��:J�ca�y�f\Jb���&S��V�s���
$)�����|K��%H�f�:��5�,M�`�*%c�0��!=r�����x
@�A��mo\A��00L*)��	��G�,I	��&��c�w�&)�y��N���
G�@�(6���2C��`�;�Q��ᐫ�� �p���MI߇9@U0�6��S%�b57�.��Au�YIhf�U$i,O�S��g�zfni0>���h^��)7,
���7�\[^G2���٘�j0hW�v�&b�H�
Ԯu`