BZh91AY&SY	<�� {߀Py���������`?<F� �(ѐ��S�G����4� hɓ@�a2d�b`ɂd ф``8ɓ&# &L �# C �ȁ�I=OHci#�d��@ �8ɓ&# &L �# C T��L�h�	?Bja�`bj~���XD+��H��T����~J��C�hcQ.*H����7�W����AaPy�L�P�l4��g�Ϗg.�ֹ�<�KYg�Yvl͖�ͱ�f�(���_��ļJ�,�HJhI.<yW,ۣ�n����o�Uq�?�2�{%2^�U��nśe_-�g�ÎwV��(�o���եk��I����8�#�M{����}��~R�=���=�(*QC#���ڄ�-yD�徰{Ui�*:)\�U�bmiv�S����Q9�Lb-�X_��	8�)չ���p-X�*�㽊pAaR�C�F��Q�'C��������5��sM:n�pƭ��Ðɱ���E�.�7/YZ��['Ưt$#I�v�̫�M	!���AzP_b5X��ZѡU�N0-�AKe��l�m5*�0ص�.��	�Wp�bp����RI��TX���Ʋ�|d�$9�iͷ�/Tɺ��v��Hx�<��Ą$!.)$��@���yC�1�cNY 
��#�#uk$�YH�i��ˠ�D4I��be!�� �dJjf�!��a�ejbBAQ�tt�tz����9��gv����(Џ|?��=�&Ꚋ��=)#4�0T�
��=�J,��;z<� ��IEMH&X�^��P�\˦Ƚh���Ǿw�g���y���P?�б���ש�n���ܲ�ix���0�\|n�jk�$��&q��H>�xG
v>%;hvO~Q/�S����jYg��|���&��m��FP�{�t
҇����*0
`����%�"/*l��]����<v�YO��9���UJB���v����ׯ����t��އ�~?���E��@�lT7bC��]�+�� �r	]�#ғ9{ֽ̦ώ}�M�����ۣn��Abų��ߎ8��늍'ED�����&>U|�GVǌ�ђ�i1P�y�@���.ҷ*�Ĩ��x`0����B�+]��������A7GP�
��PZ������Zͽ}���%u]�g2^)���r�������qn,;�Vpu��h�^Sz�S��2]Zݣ0�����u�"���5�yf��M\��0fR�V�<T�JF-t^���&�V�ԧ�z&6�w�k�W2_�|����`[.�YT�n����MѶZrds�m�Ć0 e�N- �h&9N�+�D�գ�IDz�x���]s&sc,訳�e�wfک�r�e��rYҨpQQ6f������"�(H�V� 