BZh91AY&SY�US, _�Px���������P�p� f4h	MJoU=4�G��P@  �F����a2dɑ��4�# C �� �B��j��~�� ��`LM&L�LM2100IBi�M#F��d� ��d�D��ZH�d����W���Uv���heQ.���{��Ud�`�Ҩ���@��Q247l2��8�p��ί���]��,�t��?/_�X�V����T'�Ȓ[�u)�^.�ԦQ+�����^n�����XE�Nm�jpބmr�v�]]P�5+X��l�[+$�L����&f���aޒIg��/�~���T;�������ǣ�!�m�S�&;d��Pd�yb:�_�Bl��9$V �ۭ���5]��
R��4"�#| =�fa-2���r�.�yl�v
c	�v��KԐ�Bd0E OB�	bcA��b+\ظH��Stna&b��޶�2�3f��e����	�]�ޓk�x��S\��]o���Ȅ`�+����qҮ�WS}����ٗ�uѓs��-��M���:А��%�$�P(c<<�o��t�r�U~���
VdT�b��"_��*PD�D��n�hDPj�Gy�Aj@�fI	G3e؈�!(ҏS�R�~��t1~��G�H:g<}j������k���De�HU8OE��GiP�M��{�(̝��t�BF���b���E�B}g.�O�y~����y�h�(O�,l9���n�ܘ���=��>\�����v�RO�����>1�N���U���%-NOo��Y�g�$�|K�z6L�J�D���t3��}-�۪�u1%1G]'~TE;Pi��&����m�LG�̹�3�C�J[k{y���\�h����t42m��̗�g���l����޼�yGo�/Q��S��0�{�0�[��;a
ZCT��?�Wb
s8n��N�¢X�nf�|ljVܲ����*5�z�n˨Og����j�7�j~�C�kKDС����a�q��������Hk0Iˮ�*��llj�:�%�3V2a����D����E��Q+F�<N�`)��s�u#�fg�c�����l���#�lzpW�ܨ�˱��3^��a*;
Q���M����4�v�mbxq5�*�j�:�Ժ�1�EՂ�Nh���ɡNs֙Z2�9jF�,�͆F��W[2j��Z��泙R����F���xX�i�]�(�v��%��Fϕq��)'�g���i���f�52���gW+�|�Γe-g�/�+D	�����rE8P��US,