BZh91AY&SY��� V߀Px���������`?؆� � J����Ɉ ��  L ���ц��1�d�M�`LM&L�LM2100	L�������4���=@  ��A�ɓ&F�L�LD�&�h&���i&G��FhjyL��@� �!* J�$@���>��%�
ZH& &���m�|�A����ړm� 2?>ӆ����8ƈ�t\��5rd�NK)9S�)��B���64�x�׀��GeHIpT��lR�|��̂^ ��=�C�=�*2�F�αvB��a%x���7(���yl��iw��� ��I��V©������*[�����i�GӴ7�pb6g���n�!s�e)R�r��sk��cvVIUG����}�Rj~�FV&M��h���3V,9�h��P"�L�a�a��j0(��j�/,�D��Pd�@`DCJ����4��͋r�<+ 
���[a�SY�7��\��CD4�#)�U���
�Լ�xyAD��M��d��"`��B��N��楌D
�toD�*Ψ�	)ց�����#��%YW\�	���*�3i&���
�2�
+!	Qh�'�5D�$!-I%����]��1�ƮM���/DӢĩW���IK���$���Q(��H�.F1<��j�$h�Ñ�M�t�;(�KH�I! ���f�j�! �H3G+�R����W�j�f���Tat$��8t���AP���.ldP�rxg�����-�������f���9�c��3޺����X@��8j����G�;��@?�)�~�N]"�{����^YAc�}�Y�%��
��D�43Q�@�������}m	����J���A�Y֒y��l�*��-�ZNW`ݐ�Ő��:�&PA�ѽ08�5tR��Q���5ʇ>�%��#:ƚI��4��R��Bг�?A� ���kE�*���.���ƚt�@q�l$��#�Q˦�����1�))�b�1�Qk���g e�W���q��P��u�SB�����Pe�y�؆��xA	$c]���� �į!���.:CE儺(4{B���nz'(�M ��8(!C��llj��o\5�䌎��9̩4CEBҠ�&Ȁ��� vmBx�H������ހ�&@�)�Z�����:����1N��B�A����i$��C8��y��װ@`3����u�H�1�f
��(������U�$8ʅ�ln*3V�׊�����u�,'P���v���2L�0e�J��d��Y`�r)+��D3�j�6���y��Ľ�>sHd`b
E�3e�P�Il�߶���6*Yo��A���d�s�����)�ߘ