BZh91AY&SY�X77 �߀Px���������`�<�<w�� 5Q��M20���L�2i���42	S	�( @ 4h   ��T�Q����4 � �� 		F�" f��h��  ��& �4d40	�10T�hOI��	�O*z��4��`l��)�|H��B�@�I&R�W���*��C�r�/K�����U���%ƅ�̘D����:$ 2�.�p�;�+t�}��ò��������e���4c��gT��ʃ���2W��!"�$kհ�8��a��>om6d3~��;��0�l�RXE�3���9vZ�c"̪`�K8r�,�v�2m�b���J�}�I12I���R�߯L����~��sՆA�6�(9@a2,�zyCŽ���_u��Q�������I �4�S��T��M�J�ӡ2���b��L�3��R�ރTD�Բ�y�[Q�eLr�d3D�f��ō��֌#E�F�T�x������2�1 u������ڔ��	&�er�c8�ȑ�H��M3�I������
ȭ�Sa��faٌNTXHliWnC��f�A�M)��]�%vA�k�.�F))L�ݣ*���$q$�*������	d;[ɫ�21!C���T%�SDFYk(KiovݙT�vDL��;&�LD+n763.4��Ue؂L�f7����bb���L�����lc{���C@�C�����%���T) x���a��#M�E$Q�2G�DTBX��56���Tle�(L�1�
�8�a��쀆QA@�5�j�D&��&ѩ�Mt���9s��<���ְ	9��;������q$�<� }� C�v��=��Es���]��pL��f`"!�v���s��E��/��/Z�{8�O��m�<H��P��Z:�M\��vt�������O����)�9'�Ę���|�Jq|p0Jr��|.�D�����z�e��/T��`]�9jâ
�R/>m�,�KF��UL$)�GUI�*���������T���\vEYO�{St����T�Vу����Я`�+��&����������4�P�ێ��tu�n�~�Wk�b�Tc~8W�#	�7K����vy��;�8׶p�,X����f�1�^H��7TD�ǐ����Gk:�5G�Ɲ�s��C��sc�a�Ҝ�Y�k��y�������BB0G��*��c:�5*�د�Tbzآ-}(�{��uD�=?ˈ�K��f��A.R>w}���G7Aa��g'S�����+�oTJa��;�B+�7HTw������#ys	
|���=���O>��T��N��.R�­*٢l�n�*q�׵1�c�ל�y\�~%��ןc��K-N�ٴةhr`u�կR�,�!�av����F������ιh�RTG�gw���C��̜flH�賟U�Vʩ�s�e�����^׎�?���)�B���