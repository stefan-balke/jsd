BZh91AY&SY���� 5߀Px����������PX�3i�uP�M�I�FSڧ�&�����4 h�����hh     !")�<�OQ�OSFG���  ��0L@0	�h�h`ba"���1&J~�5?Sқ)� ��Q�3@=hH��@b� ���{�Fq�(1`РЬ
(S_��v�=�,�B�f,"h��4�#�vM<5�8]����#� ���}��:`8�C4FĲ��$��)H��v� ���jQD	����U�HԜ�(38���Az��:I )�t�$
�T������H�"�G=�����گP&6�M���iu�r���K)����q��>�ƕn_�f����,��6f�{24��#���'0��Y�HpQ��HyMvu�h��!j�̑p�,c���iQMLvZ��F1S�@�<X�cb��j�����t y�)��`�㋰�8�؉-�S�gA�o3m��Сk��v�9P�;�j%J$�f�:0���q�X�6If6
�1�����V�)B��PP0s-rf�`L¸�g~�:�m��E�`oV�ǌx���!��Z���~��e�"'�P��{�5V��j��6T�bp�0>�=V{fDs6�}a�ɂ�M���B��J�����8��Q�v{nA ��=B�}K�f{�\�� ��b���҉T�n`Iv$HcPfG��͐ |�9$���iK([B�i�h���K�yk[W..ŭ�B��0ka���*ć��D�pC�����w �CI�a3�aP�!��>�t��f�1`H*bO�xw�L���0[6\����E�R4�� լ�X���CE���s����Ԗ� �^x��ҹl��oY�� �זa�{)JcѢ�X�'o@.�G08������Ӭ/*Cy����&JD�aH�Ld�"�� 
8��"���萍/Y.�p��7�"79�Ԙ��P�*%	2_�ݹ	�<�z
@3�#����=��� 7{ fn9����c�����;���'��^|���-jҧa�,"���m��w@�z� 3Pm�ӑ�i��f4�ሩR����X�"D�
NۺI��tF@�4yx^5I��Å-��F.�h�z�QiH����t�C���fI�s1l��փAD����X�7� ���m|��u��Xk0"�!�B�����)�E�%�