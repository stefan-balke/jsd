BZh91AY&SY͊EJ �_�Px���������P�pn�ps��� 	D������3Jz��4�4�@  �"D @     				�<�~�j�m  �MC�c�A�ɓ&F�L�LRB�A�SLP�ʏM'��224����bH�r�P�"K!_���[a���K�B����Uc�kR@̘D4wZ�Q�	H�����ϻ���y�;��lh�Je��7\���H+x��6�w���N�(�(��>n՗5��0dm�Ny�kOE:�=&�|���tF���x�I�a!`2A�C��C�Z��(��b�/aEUE���gr�<H�y�VV��Yp� ˧��P:? �E�@�.#OCvR^�6+�t�����Y����H��P���ު�`ZŒ���JT8�i2L�(C=^a(�s6��"D�]"cH��VA�\��d��E�R�C��"�E�gB��+k3�D��b$�׵��X$l�iV�=(��7F+fdEߐ썌lc{[m���B����*K��G*��w�(�_ �ڒ6`]N�T�Y,�Ix7C�!AZ"�]�\e]"�E��$Ɓ��][*��z��V<���g��끃����x�7�a�)(���Y1��0Ѫ{w^K�%���-��f��2#����c�rC�����w<��?���荞�!��B�I���-�q��0{�Z�?�����4�|����5>Q_�f~J�9�g�LJ&Fr�G���Q�i&��+�W"��z����Ѽ��+".W�a��e��g���Ss���i}W�~������S���aE*%[����B��y��u���t��L�ǳF<�a��YuuJ)��W�E�ל}=��f��S;3������V����֓��a�a�So��>ɣL
�#�������I��.9e��>QRn��I:�懿��EG�?b�*��������5��ä��X��{:
;[�Ab��$$#�%��d�����M�3b-Q��glR�-���:^�ؕl���|�ѐ���zK�;�4>��MŇ���w���=��:Z�#�Q)���z�����%(���!�'˄����Ƴ�5>�͆J�X�;��X�ʭU��V�3S��=���=�=���K�c3��gs$3V˯eZ�M�iЩhrdsɫ^��4T>�W��^_8X�/����u�{�IR><<]f���Gf)��8^,��c�ͪ�~nٖ���84Zj*&��My�w$S�	ؤT�