BZh91AY&SY5�&+ �_�Px���������P�x�c�i����?!=SyQ�E4h z����ɠ���O�S�M���@       �SJz���dɑ�@4  M�	���dɓ#	�i�F& �"A24&)�4���Q��ѣM��l���"$�$�� ���9�C�e.��6�CH�Ms��ۂֱ#A�f364q5U"9G��7w5v���f�V:��''S�m��-K@��ʡ���X��������]�*2�F�"��/O�c��G��`�x�K��HE���0P�?�S��rqO��<~E�0c�W��x�B.V�Txq�d�i��.[�T��V�/�6;�)�`�Ɖ��J'��U�
����sV1��<�!V�[�`��U_D�B���Ū��핬��$J��G�B4"5�u��5����uN4$J�[m!��7{�㤼��x*�Ë*�����	��2yIs*U �ci�wY]@҈^�A@�5��λ�DT4.��'�j�lE��T��ǎ83��h�,X�j�f�!ՈͲX849�
��|gj�A���jS:z �{�C�a�A�W�.�x��o!��� ��3߰՛P��d.c�_<ᯭy�rKϼ�^ y�K6��gSb�,JcP̊���A�,�z(�l��7l���1cPd�E	v_��2��0�Р�0k^e��W7�a��36V��i��LbS�A`W����=�\k%�*���.��x��]Z�\�Y%�I*��U�B�{ɑ�6X�Q3�RI�X�VS��� �/� ��QV�ȁ��[Dg^z�0�ֵ��چ��e^�<{�Xe{��l2�^rp,%�*00,6Z.Θb7{WSQi#b�(,�	�,���$�# �+��wf	�*AQ6Dfۉ��BySP���c�rP0AF�]@u��x,<�H�E��t��CBe8�� ���h�a���1	��x��NӸ�8��ʅ�A�恜8�Ɗ8D�/m���f[7Z*�+xn��n�E��Rw_��/���dhZ8� �@�K.��Y`ð��b䪁��c/j�F�������b��q�d05�e�Ř�d�7o��������
Yo��N�l4+�.��.�p� kZLV