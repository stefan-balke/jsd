BZh91AY&SY��F X߀Py����������`�<�` 8k�@��U=�)��ѡ��F�   ��ɤ��hM    �  sL��Lф�hшd�� A)�(��4�� j���    sL��Lф�hшd�� A"!S���jz��l��� ���&r� �H� U"�  @������ � �B�`��	2Z���8?PPi+ L��SF֮�!!EH^�񳩯zk���'c��2w�c��󙹷��6�����t�t���\�D�y_����zl]�J���Hۦ��8�H��±hƱD^K&�Ù���
)��S���=�xhх��b:c�gOA��
*S��j��9na�-E6a����0Z����B�i�Z�Ap\xdo@��#ah�dϛ��8鵭kX��kF��xB�|�]��l��DTPQg�ҸC�Cib�-����*�ءIP�R�R��"�*~����p�}v4���dt�Gr!�z���<�I�!��Ԛ�kL��jS����PP��K��F�f��G5��Z�o��)�v�ͅ���f�����%f.8���B�����[O�4�d��S�N?B��#�lq�>���..L-�u3B-�3f��=�z��'�wlכ�W+R:ڌDL(�˦ӆ�YZ4�lӤ.r�}m�ƌ��re�uޝ!5���!�ÝR뢤�&4����IC�*Jփ/[M����fU��=��������V�٫��F�y�.���94
�q(m+��E9A�����3@��:Mz{8�QpEJ'��V˷�GDs;=��h�����=�kS��CDqigN׻�*�Y%
x��JWN:+&{9&�(�"��U�
��6�c�+wp�*�f�%�$��iE�DR�C(G�&,�D�`�XJ����X��ZK#*�D2)\�Q�LIAK�$$�t�'9��F��5#ê���n4e�>�F,���r���r̤DOqq١
����)�,�M=7���L,�G\���2*��A��s*��33J��(3��.=����I���-F�Iw9�wZ���=��W�B_�B!��r�ׯ>�~���( r�eBT�Ҽlޒ�P	��!/�0f�¡T����w�Q4�C56_��A�/�I=5	��Ʌ��{B^C��3w5�B$��9g{VBL����oM	2x`�H��M����6̇=�%慓΁@� 8��p�����|�5�%�QHX���;?z�LTHK���.D�M���-�{� *k�3R�K��K�B9-_&����쒼�"�/�jbJ�>+�Xf6���lC���'2B]�c��zG����C���!T`h(g�$�I�Z��<�A� 	8`�D�n��!�/��	�E�(MɌ�_#t����Z,��$���Ϸ�j�_��!.G @��04�G���xz��J .�9���m���Q��hL���8�ĂK1P0�3h:���;
BL��e/9c t
�{Ma�ꁜ��$cB�q�Re�q�!a�8����خ�����pY4г�q�a��@�(f&s8f�K[ʇ�.$.�hK�u��q*�@©T#�>��������h� ���#A�	Iq�e,$�� ݮۻ3k�ګu���h5\�����)� ��0