BZh91AY&SYԳF� 7߀Px���������P>t* � J$�Dhb�bb0����i�M1�	���dɓ#	�i�F& �)���MM P   sbh0�2d��`�i���!�H�A4�I��&���L � x�O)���BD$
�bH����# AV�!�LI���ѷ�A
ᤙ����6�#�����=�j8��d)f�2Dwe��7��
a'm����b���x}y��Q��>x�1	��C9('1e�wY����;&����1�y���ȑ �q"^2����-V��M0cۗϤ>>�F�����k�%�^,U&�UG�=������f�/h���<��Њ���%4@��EH�rf�j��s���E��dw"�s�,����1V��ű�g�����������I!fb�j�e��F���I��i@��5����dѼ�	HBZ�I%���d����1�Ɯ�HV}���.%�M��b��L���sx$�r!��a�a�y$$5�V�
*���X^U왒���֧�C��(F4=�O��G�S���͸뇇��G�X"`T�T��ER��Yr*�1�1.�y"UW
*�b�*	0;����83�ĭ�0_�Bă�0:�i��a����4��瀲⾣,�IyrU ��G5�#ơQ3kb�X��!���k ����I�J���%X�b���f,jl�P�M�	��nM �&H�T�)L��\�p3��,3��p!�8�P�b{� �]���1q�PP�b)�=�����)��CPA�!z�#}Q�鮀�_A2uCE%4-o�;
,�:��&n_�~A��n:�3��_%�J3/,B��k�ْ6
Hд�]�É���zG��k�^qZ	mG���4�)��0Ү
���"5�m�A!C��llj#�;D7GLFU�PJ���(%c�n�y۵	�0.�r��{t$f&@�9����� �=�>��HiT�r#y�m
B~�,��0�ِ-!1PT<���OI�\�o��A��4tt��Q�$8�Y�Fң1�n�"����sm�,'P�������_""�0��jl(h[u��E�\J�<T��X�;F�7L�M&ă����R,5͗�KT��x�mmx,���i1!4)`v[O�]��BCR�X