BZh91AY&SYT�nu �߀Py����������P:n1� �QM��)��OM#C@�=@3Pz� 4���L���  � �    4�
���hz@� h��   ��!�	�4ѣ4ɑ� �D�L�@'�6���4�  �'��L�� T @����r3��*Ф1Hd�����p/l�+��a�a�I�h�������R�tc��}�w���o���a�a�d�A%�pͬj���b�p�r<Y��H��7�.RFD�"�6��+IWc1�ރ��y&	"�au( ����#��|g��9,jn�
*�(��ʻ��B�c�	���"��3e�F
����LaR+�m%��ޢF�u
Q��C��5`�0̆�4
���[�S
Yjb�rb$�Ԃb�6P�$��$%HE�Y�Y���X9�������w���Rbs���Am�k��e�A�	�$�L ������b66�)���n0�a)ȟ�7B�(مPpLQH��"H��F$��1&��hJ��`�)�UATH�D�_�`�v�)u�IT��@�<z|��}��p�}��8RY�H�C���<��5I�IYy����+/'�C�Â�����Ь#��� ��2�o�};3k�T7�$�Ā�W�eM���͜R^���kؑ�͇�����{�i1��j<�G{ ��d�I<(�r]C������A�����|�5D�#zg��]5|R��X�gEr������]ވ�������� {n��*b���O������zH�顱���$�VGW:��g��-�F��tB���آ�)���P�e��hf�ף9�#�ٖ��^[(�V��~�03�) -;�<;N�:Ju���U�g,F�A���\f��B���!
�G,T�L�����}�AD��:�iX���PRh�z�!D��n<��=Tґ�p��f�y��v��浙Tͧn����j+�wā^G 0MA�9ԋ��,UŎg�d�d�P�0Tm: g�v���RE�`�%Fl��V[Í��2�MIߗ�D����"��P�3@���Ʒ_bAku7Ia��P4c���0�{�4��>r=F���֤X֯*Io{��}[�6����-k�Fhc�vr��H�

�mΠ