BZh91AY&SY䂎 �߀Pxg���������`�zl���   P	���#�L	�   ��dF��C@ C@ L��42 d�  � ��Jhd�<���M  �2i�# `F&��4� �RBBi�@F��&H�542F�m�I
�-&P�H�d+���_���������K�	��L�f*��0UD�)�%G���Z�Y$��"`�W���-��%�Ӵ��L��3@TQ$�9��3�@�oQ��"ًp��1�K�25űi%>9]��W_���ݮ��c���۷,�+V��h���A�Vtq�#�q����k�]r�&���C�'"Ţ��x��U{����hk���Ϗ�������E+�n9���g~�����+.D�S�cD "*P�NbS{�%����050��f
�[��;5��.�4���|�X�V��jH��om�m��E�E)�v���ml��3J�f�mg�j�j��Cvr�Q@I�MBJ!ô-f�Œ��cm��ھ/l�Zi�0�f���l��kj�uتҚ�SZ���v�4i�"j�]����
8��*����Uȅ ���&P*�I��2 �E	������t44"�R ę���� �(�p���O��U,+A!` 9rI�-́wd�f��Nv [��	DĊ�!�!�;B%��JH���!G	�%�*���Z�z)�/{ܖc[�%2BL:�
���'����?z(¡JHd�3@�p��\��
 ('T�h�N�P���`k����Ҫĥ{Ib�T��T��kl/���<)����������XSo;- �'��w�{>��-��6t��-�]z�S�Fi���8\~S�\���Sgt����8�؃��4u�9%;huφ�J�KS�#����=�=�J�����f�s��R�V�Sѻ�V��r��%��m�S()��y%H��M�K祦4-�O3�u>f�_TYU��;��=*�{��wu�Z+W�X�S�?��˫�QH<�:מ���8�x�����as�qQ��2�ν|�NÄ��a�M�.��ų��4z':Bŋo��3r��~��Ȩ��:jIϵ��Q�g�+�Tr���</ܓ5�0�gj�t����qab�/d\��-�v��Z�R�k2���LgN�3���ٱ���Y��)k���OglJ��3��x!N��E�G��^�����,<��ηs�=��/V�9*'b�<_3�l^A��⎨*8����Q�0��MZ=Ka�M��5o3T�YB�
]JFuh���I�������߽3�g���N��a�-Kֻ| ͭ�,ro�.�z������ٷU�4TvW�t��p���7���Ԏ*���RT��g���֑��tM���Y��c�ݺ�wl�M��*�%]�^̿���)�$p0