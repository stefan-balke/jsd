BZh91AY&SY�'�� l߀Px���������P~s�utj� �E0����!�3P1� �A��S�#i��� @� ����T�Cj0���щ�224h�9�14L�2da0M4����$�4�$4&51� &&�5�\`��I���D���~j��+KJL�ZT%T����U�}�M*��%�H0y����/�[�{��n���p�:�gy��s�Q=�~�q���� .̗4������@~�ӿK�� ����ƫ]Dhչ���[�u���l��Ucy1ѳF8�3=��F�OM^Q�����{�(�q���N4�[�#tmǿ\Q$Z�AP�t����73��M��!��1����N�]��sQ���eӶ�3S=�-���S}L��X�a�
�E����16�0�І���&-|�>L����kE�c(1u�i!�E�X����vJ��&����k4׫��Bܰ�q�$ÒK	�>F��S�(�"�UV �N)��<uˉ,Ԕi�jh�-Mн�$�,]2�2�7���Г0�E-��ZXKT�]�Eƣ3ta�$�)u��f�C��R8���"��8�Z|���*�8�Kp�U���G}�3\s���j�D�;�+�,�r�1`:����9�0�^�d�?�}�d4x��б���W�ϯ�.zJ9�R��
q/������!`�L�E��\�FXGr��p�21R������h�s�3�HZ����qgyޓ#��bKp�r���(�r�%��\����i�Rݴ��*�|zٶ�>U�I*���]f^Ev��w4�9�i�v.f������?<��ǁ�=p�D�v:o��*aC"�B��SQ�&�z�r)�緫���h����Z��-�xk*c]�(q�%�*���Qa ͌�
�/�U��&���qL�7.m�R�sZ���ۗ�Mr���4�03b�Uu"BBvh����Z���<AD0�2=���k��U;�ǟ�J�@}�⛞��3]d|���v�wV������+�{͂���Q)�[��f�
���u�Q��wCyqw��if���������Xj7w���C���4i�	�M��6&V���u�s����W��|�mx)e���n����M�%�Lά�z����6��B����T��u�q��ԔM�c����v�L���E���{�l���z?�s*TM;�1��ܑN$=	�� 