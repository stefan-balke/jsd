BZh91AY&SY���� L_�Px���������P>rl
$����L�I�ba� @h����M@ �i�   %2MOPd�� �   9�14L�2da0M4����$H4d56POT�<�LG���4�CԼ�@�I"%D �����#b_� �HSd5�/�m�<f	jɖaDm�
`[`X�_���߆��/
׶���@'�@x�|�h��lW�&�uT��;�N�'�luy?Ař��"�,j1�/$lN�l�St�4����}�6��c�1 Wl�](�+��g�ظ��W�I�C�̘j�������i�nAu
*���j��H��SBFX��b��jN,��e�� �@@*�*e"$Ce�����HHz�$ь$���a�%"Tv��H���(U9E���*]u�DB ��fC�i�=F�h��U;�:P�)6'K����r�"���VdǄ�"B��$�!Xcs`_�~	�@ӆ �'�Àܫ2)��S�H6��LL��(�XceZG�ʌ��5H ��	k潛؄JQ�p�_�͊��Q����Xnb	w��{X��qC�$�z)�8s�P<�|�4�%���o�I�Cn�&L�An1�3�b�;8j�8�rK�&�Lk/P~�`g�#	{�8&	��Z�Р@ÐKP��D����*Ғݚ&���"����,������g�w�� �-ڒ{h�n��J��Yf���E	r�5D�M]	��0k\R��R<�[��g�"�ի��J����� y��[��WȠ�'�;���Sv���v�2	.�H�9r��.�Bd*��Jh\w%0mS<	� �~{zy����ٔ�J�r�����A��Y)�C"U�H\4-�������X����8%��00&X��+��0&�� 	[��L�ұ2 �!��"�A�'ff2e�D�D4X=�@"l�ٞ����ȮB]�@P`{0!��}����mĘ��9���Bx��>��4&S��:BĒM}0��ԉL��d��<0	���A�恝=�*8D����3*3~Y�a���v�bu	�%��TJ����ض�P����ڮ$\4��Kl* a�u)z�Fo�3I���=��S$�X�k*2D���{k�f�k�v`bB	�B�S-h�ܑN$;2�:@