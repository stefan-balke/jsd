BZh91AY&SY�p�+ �߀Px����������P�97nb5��	@��)�)�mF�H��f�4�i�h6����   �   	L�e0���3Q��M�  h�& �4d40	�10� SD�	�)���!='�  =Ѡ���	
�P, @������I� �B�h	��_��n�4��hVL�I��R��I��-��8qƏ���,��̗Lyf�(�������r�b�Ă�y�5"J�Y&�i[�ܯަosg ~���a.2�3�hO#�A��q��i����4��z3�HU �zA��fŸe�IW7�l����q!0c����4��Y�)p)Y�a���*�����.�����d���q��V�e
]�D<XL�QH*#(�U��&�eb꣋5ҼS9�R��J,g����3�:$�vR�<f�	��M)�{��bZRt�j�*1�C�����7��A�;�
fy�´��*@j�(��&)$��7
��T�L-���kV�;�!ؘ��SE�����uD�$!-i$���F�0ߒ9xƜ�H�G.F���z��آ��6�m!w��YX8���T��bW�B �y�� ���/(���uQ�UM�鼴�k	÷gw~��Νd��z��5���Ĩ���BQ.�m�N�����JY�-F'��-*�hJ��"���t�;���H�@Ў���#��8ـ� 2 պB&ǅc�I|�Q$x!?�`�G�aR��d04�|����|�]�37zI�@�k��V���t���Gf���DP��-�PC(�����K�C�M��L��x����gÑcw4@� �"�A`�� {.����b�(
��<��S)�Åldפ�7����C^�D�����ݫaE�/S]Ǹ��-�e
�?�Xd���ՋH�8�/�!�E�nHb�aH;P������q+���UC9�#r
	��"s3���1��!��a&�|2	
��
FƢQHe���ih���PRh�|�DM��BY��ՙ	�=�G�Δ�2�Ĕ�����f,j�@~k6�Ķ(f&�鏐j-���abBC�"3�3qy�b�TDϖK9c��>���+�X3�MQ7�!�c��1�#��Pf���a�7��߼�*�Q+� ��R�f�M1���T7Ե�$��v�Ib�XMY	����K�H��{15��/"�F����"E�k9T�$��:�@}]Z^f�KZ�͘���B�ү���)��iX