BZh91AY&SY��� m_�Px����������P��@i��&�$�m�)���h23S�4�h   � �`�2��JdBi4��OI�55����5=@ ���9�#� �&���0F&
�I�S�$ވD��G�♨�@��2mO#DEtA-$��!��d+������=���DE "Tx�$��DFE`F8�b��mA�~�ǫ��.�1���^�=��c�(����[G�yU�+����	)|/R��l��.�GJ<[���0I��[\�kz�2eK��i�l2����h�+����~�/�	�e��O��;��nz~lG0$���c���ѡ/��(]��M]+(D�c���u���+E�K�V����r�g���"�t���J��(/���i�������	�5��{����Rf)"�;����6�:�x��]�H���,35RB��S"��	�/>�0n�bt���2H���;�)2l�o����e���k�y�N"B���I@�3�GO`uI��NY +?D�\��j��J)M�J�%䖉s��Ƅ�.j�<谢��3+HH j9F�BB@%��be�S��������@LDD�;_���d�@8�]��lJ4�NF|G [�e�{wZ�a�ޘ���%�ٙ�3a�#:DddE^D���9�39�hN��aR8��,m6:���g*^p)hX���4o�Or���>X����o��vS��sیMjf�`}��Yg�NRJ�yvi�{ti���U�K9ih��:��x���qPC'�st�&L󣮶�1�WidQ*܋�f&���ҹ�nkzT�\��%�֕�3��{/���,Pq�{�)�e F(���
0�SALHd\��X�0��M�D�d��)������c�&M��ղgP�V�_���l=tp�S=�I� 3TVGJ��vU�9o5��1[<�(d��P�8U�KBb"5$���V�
FƠ>�� �d&��bUQ^�ȥN��-���m�ܑ�|��+~�S�6��eH��������(�t�g���Eѹ��]Fj�Lx��s�WH�%F��(����ƅ�驥��j:SWZ�R��<��)�n��B�F�kt/S>Ȼ��:��qĘ*�Q+:� ���cA�ll��Q�,nX�,��4�;�L���@țR��H�������a����s���6�9���_��x9�t���Ȩf��kɧ�rE8P����