BZh91AY&SY�أ� �߀Px���������P�n��4��	I�z��x�3	�)�bdhтa �S��� ��     S�Q�E4�M@=@  4 ���a2dɑ��4�# C �!�
m�ة�ڡ�?SPM��꞉��`h$@���H����G#B_(ASB�H�C$י�6���,�B�el	!e�)) �E7	�"����4�M� ��J'����<3h��0���Ek�j��I��z�S5ePVf0��4'qIH�����T�xO���S��4$�.�=( ���?�Yc���+�)m�;4��Cǜ#2�Zc�I��>��jR]:�(�v'��u����"�d:[n�f���fɉ��oW���cfY���&5�t/|I�%�C*��Mnش]1.d��x��*�e�����M#�E����(����!I��^@��F�"Y�(g�D��ƪ���.�&7�a�710)$0Y���fe* �	�HgD�eTK}S��,B��r�&��|y[q���_�iՐ*��Y����x
)�;��r>�E CIr�)>6�¬�`,�b�)y�½IƊ	�'�[�{@o]!�sD=�P8������h�����l�4�_��I|�EIx$|у2>T
	��/:�6�62�e��� �WܒwP%UVYK� +:���Ơ��E	p�6�@e�3�� ��5�)T)U��U�2'爹�3�aTQ!���\-�;����%�
b��*'��w�4���.�H�R8p��,�i22��в^�e�z4�P ��f�GIe䨅=%b

o�-5UW-���r����+ڑ��� h�+���e@��0���Ш`^L.h��B�nxNQy1
�Gf*H&@�TL�"h�I�E0w��6�t�Y4CEa�T�d@F����P�Yd��n(/</A!��Kư�/5�%� 7�n�����>��)�����@�`&� ��kH�&9�����+8��i�7u� (�g!
b\ I��`�$�9� s`,���8@(,iC+)�6G�6TL�o㞙�����0Ė2�K��\_�z�54��>�F��;PH�Գ�#"�`<����ة]��^`B#���٩���"�(H@lQ��