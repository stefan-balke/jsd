BZh91AY&SY�� ߀Px���������P>r*P�@���I%2d�5��d�14  �sbh0�2d��`�i���!�Jz��)���H4�z�  ����&L�20�&�db``$$�L�����=5C& h�mCSF$�O4�B(�,/�����~×Bm� �B�b�1�Q�p�\��`�a1BF6*�X� 1���͛�p�c�Ӈc �;RQ?~���\����Ɔ�"�4iyN����H�R�S]�#��/Nd9JB6T��F����$���9�CR�ٌ�\|���MpV���2��!�wa��]�q�N�:V�{(�fM����Ļa����9�����x*�%�a f	�qb!��cTP�L	�k�D���Z.qNE*���d��nb0�R`� �i�?U5��M�NG�3
Τ�xh���8�EE��5�"��U��$���u�Ê�7�%���o<�MM6�k�6V��*eD&���&%�Ģ%�����!�[:((�7iNCJ<�i�y��L�>l�p�<���|4X�r�O�;�J}Kd'�Pf63�x��W���Ǐ�u���1S�t�mS�	AU�q�zC��a�R�#P9��d�n2囂�/V�	��N��/���jIk�H�L_`��53a�@�����_�C:����� �]D��J���Ɏ�E�gv�[��62B]�����P�δ�v�5�R��R=l�\P�gǰ�Я� C�E��^#������%1@P�^�?Our�; ��k$��#uQÅ}v����vCEe,)#T��Fr"�16�0R�����&�A��p:u�dku��˵J'Ҝ�!%B9�P
���a����Y%��a��@��9�!hnz�(Ț�� $p�P"A2J��("b���EC �Y�e�9�&�h�zJ��� #F�K^hOd���n#����0��9�7J�EC��a�qI���?8k)�w��Ē��4v�p��# �&|�W�;�%��+���i�7n!�ST�"c��\fTf�����E��4��E��&���qA0��q&��1�`��*Կ��4w�𨁄+V�r(��C�5//2L�!�Eа�A�)��)"����ک�ګuJ�Ȅ�
:�#�rE8P���