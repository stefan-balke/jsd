BZh91AY&SY��� �_�Px���������`C��\�  ���O�6�= 4h�i� �0&&�	�&L�&	�����Sj��h�� L�   ��B( hh     �A�ɓ&F�L�LDB&�����=1COS�F�@f����M%!�BUHJ� @�?��rj@/� �B��T��O�p/J��\�s@4x52C"J���7�ye�n/A�.����ӭSM'GGQ��pRQ?~o����8�^6��%�EZn�\q�DA��5��w3s7m���\A�tv�A&	� 22ȭ`ѕ�1[�J!$���$�@~��i0g��.�F�F���u�L�A���OO�P�m�;������^-��:�6��,�TeK*YK����!��)!i�	h�D)V���Ѿ�%�%#�a�递����3��%ZH��6�n����	4֖6,��w�R&2Lh����ɖ�b�Z�/b�.BI�Q:,S$����M��7��R���T�b
��Ɉ3B%�Vėe�&����d�D���o���Gs4IhHdwR\T:����@��C���D<��DcIq ��ɴ�(����%4,����wS�Xм,�����[FS}�7�o0l\��NO�(�"�[hhA=�Wx}r��Y$�D���L��	b� Z�!jJ-X��7(�#���e$ɚX��DD�$�I%J����h���$��k���bC!AJ%�/�����m\X~ �ѣ�S'�s�D����@6�� �I*���d#����t^�f�F�)Ca�9�����W샊���y��X{���x���|@dOn�=�N�
��BdE�H����F]�%S��҂�$� A�F�f|j703^� �`�feC��dzx$�5	���Z��b�ݚ[��6�Rz��-T@ʂ7�nM$3�E�"��6#͜�z����bƲ�.��-��@�h�6���X������͉��3%w�VGo]��~|
��E�T-��=�V��P�(u0���pj���h ���H  #R�fG�ַ��h�d���������-�>�æ����.'��"��H)C`Z�y���eR�� $�t(!B[E� ��~d�T��4f��,Q�`��"4�ؒ��!<��;�I* �O��#�;����j�(7m�$�=�>��4&W��p�B�P��:��A����T�ذ/;N�@{e���t@�\� �\"G4�%�g���Zl�	,N7IqK�r*,a$D�����(5��+��V:���A�Vp�T4���rS��25���f�yu���	.6�$%p��Kk�7���f���������ܑN$8Ad��