BZh91AY&SY�7j� w߀Py����������P��n��C�����Hjj~�hI��z����i�4ڃ#M��5=&@SԀ�4     		EA�=@i�4Ph   �2i�# `F&��4� �E4M	�����*~�j=S�i�=M dFɐ�Iz@��"�JB����`^1M
�B������n�`A�a3"h��R���4|;�����^W�ߘ��X0�5��!�0�y3�7:Ga�B��K� Ӌ�&H^6H��=���G>���q�9�	��p╈�}S5mȂ�kPЕ	$*�i�P�.��k�M^:�����g��� i��~���2q�ap��l@����6�t$�I�܊3��&��.��[���N _�4�-��ԅ��$]���c2C"��x��E��,��B� &"2$��2�*	�ҐIL�q�1a�F���8Y��W�":�J�3J2�Ò�-b�x�����	 �״�X����/PV�f���<*��c�U:�#plcc��m�4��r���и�Dr�Bw�h�(�ֻ�Sn���1+&6�#t����F8H��U!p�F]BإA@�5��; ƀf;Z��7�t��'�\58�׸.�g��⹉���/��t�F���L����[Ɂ���AZ�3��$s�;M�6�)�帊A���u�}�w@q�?�a���XD���O~^/��$�|��y��͛�\Uv�>(�dl<$X$Ά����5���-˭�$AwRI�@�,��'k��~��%#[$�P�|f����LHd}5|ȥ�\�E���L�hpg\��i�(!�9����-Ck9����H)��y'!�6�Mt�hb@b,P�c&��¨��g`k̂K]Ѣ;
!`ެ2�YB�*�%4x׀Q�2F�K�Т�8��e���=��¥U{�I+�l�}`4o)�|�H5�.8�������`Ҝ̂�7=3x�&�f�T�@�A�+������gD����.(h�>Ҡ�M���7yf�'�V��z�Xo6��J2G�/��6PZp��b$O��c:����î����"�'Y�-! ��!���04���Bb���\T�u�H�P-�(6����1�W\�-B,�e�Y����!Y$Yxgz��
��&��~��d�3# �5!CY��+n�Z�^���3*���M�#A���bli0>�F�šsA�PTد,KL"F�R�n��qΩZ��3�D`d(RO�rE8P��7j�