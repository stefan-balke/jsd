BZh91AY&SYI4`�  _�Px���������Pr"�1��40�J�i��2��I�h�i����d44`LM&L�LM2100	OQ4Қi���4 �  4��A�ɓ&F�L�LD��A4��'��H�= 4&'�yLI���B(�,�@�����r�6�U�I0S�5�/��p|��hVL�	;�R�3!���ۯ�a���t�l��%����5��#'A	ΨF	`�Ԛ����K��e�X��s�1Ă���e�m:�Y�k�ϫ�Fkc��0Ia��X(\o�$�}(W��,o(4��ퟟ ��^��Ų]�t�$n��i�7��Rb�?_�1�_��\�WT�F9�i�RX#ȅxa2�Հ�bŰ/H��67��3"��CC1EH�j���eNת'��s&�{�/e�H�e��<�2L�!P�R�lEt��I'w���Dru�f���z���f��	͌K�T���QF�]%��fd#��%�C*$�TPP!,o��20�?R�aW^6bsz�KDܔ���AC����l��у�u�f�us�q��q׼|yH��%v��Uli.�W�6��Xl��cnF�_���u�DH0 5'C�5�^����tm$-u��Ex/��r4/,J��#�ٸ��(&o`n^6B�!�P=�̂�nēʁ*�멥]Gk�q$�r�g[�.a�%(��XE+
U#����x��+��q�C�`v��`�����R��(K����MZ�#�CfВ�$�J����o�/ۼ�ڡ����ٷqE�4���@fyzw���Br"f�"�0���kyl���:P�F����v���W�}-�� �Ib[£I0Ɋs5a��9F�h$#�R�	�:V&D1{��E����8�\�*X�$� �d@E��~��Є���GA�&3=���&@�9����d��q��G\�5	��t��$��Hh�4r�q�Q<�W�9Β���*����6l�KE栰Θ3�γ6qo�U�W ߁���,N�5'~��*a%�hZ�A��P�RW�H-a��Ie
�i~
}m#/7�#�����sz�a{b$Xذ*,�7q�|x�mx��q[�����BG�����jO�w$S�	�F�