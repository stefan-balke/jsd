BZh91AY&SY�s�� B_�Px����������`?���l��T ��CF�bi����� 4 h Q(F�Q� �4�4 9�#� �&���0F&�&���M24��FF����� �`�2��H�Bh�	�!2�jjd��=M dє��=� ��B�! ~?��m�B
�)&�� �5�?��^E�B�2�G��ID������F�_]�jv;:'�hә���n��QjaBr�|�����̂�ee(IN�UcC�<���7��脾�A��{8L��H��LG7���2'��-�UE#;0a���{`�<��B@<2[)��P�`��Ϥ!?'M�)�.��|��G��b� �L��@�`wt.t��[ϻ��S*����!CD#++�9}�l���)*E���b�hEIt��Y�@#��D2�T�2�-,i3#TL=@c+Y�H:L�'�3n�.�w4<�9�%U Ya$Kb�9�3,9����tA@ĥ��|�Trb�a&! *2	�L�����)9��TTN{�FB�fa��h�X :N�	��Ĵ�,V�¬��!�jJB��+����L��we�^�'R��`<:SB3&��T�m���p���7���hh;&k�Y���$�Sޑˑ�X��XCM�@�$�G�Aa	E6�۸�E�	Q	C��1��@.�Ljr��IA:ȐHC[���llm+�r�����k�[f=z��&^3��>=n��T	��'qE�|)<���@%�!��rE�0_�����-p�̒��l�H!y[@���o3���sn��C��H���B�y����Yt����4���%逊Y�^C6r��J�G0�F,�yP(�9����L�i<��c ��-ڒxP%Z�v5m�u-��N��֠��DP�[���P[��ɡ&Kx�d�V�G��+z����RPc q�C~��+���Pg-1S	u����S���CS5�I�#����մ�a�l��T-�ٳiE�1\
.�02�L9�/з^|��~L�SH�p�y�Ǣ���!�2��;͠w����/2�����`}�
�AA��
�8Y��ĒH�� $sgP"A2K&9�9A�D���J֋\�%Ap�,6D_�6�K9�ڄ��-� uҠ��J��=;b���6,��83�6Wږc��c�Bey�i�,$�0 hy:�Bb&y�,:N���+y�e
��Dݸ� ɥ��!s�y#qQ��n�*�+�7dKu�,'P���')@�I7�6C(^5�[�z�]a ����n�͚J�0��u��=�m&�A���4�H�ԲH�H��L%��ةe���h4�L�����)�k��