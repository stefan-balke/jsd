BZh91AY&SY�Nd �_�Px���������P��Mݠ�q��l�
H4d�?�Tz&F�(��z�� �OH5=2��Q���� � MF����P��   6�0&&�	�&L�&	����I�d�54����ꍩ�` �C	�bI�%$d ���*>=���6��0Щ�&S\���p[�$�
�e�@4rjRċD�q�ӽ�����Vwg����'d��N�Z���>�?��q�cz�s�;($�E/�����L�W*��6���1�tʌ�#!Α��'��KY����&[
r�s�^3IZ��*��&�=찧���3�����~^+��d�	�k'�������G��AN>6�Ppф^�t"�m�J�ڟl �6��0Ƚ�NuE�EAy�Y	��س�Uf�U�`�QN���*,���x`�\�SU�@��p/5t ,.Q�%�y�Ɋd��ȥYv�ep�2��T#G�f�!�4���,�ˣg��٢�-昺�@�un5��I��P���7!Ƥ#�I��j��ccޖ�m��PAˉ��<rK�����(���*���*�7�8�Ld���P���wH�28BBHE*	vYc,��B�A@�5�ћXb`���g{7�n�[J��y�?f�u�/�V����a�p�<��W�7�q+;k�&���|ⴕ��,�����S0�9��x�u�6sQ�]!.,��r:��/@r~�O�0bq}��0�B�ń*�����_��lI}�a�&#ցpF�(wD"&1`(��(&Ø���d|�w$�����k��F����va�;5C!%�ͪ e�	�͉A�D��"���������5l�4�m�4'4�Z���l�ls@�^ViQ�F�͡��J�� \o
\�ѪH�rJ�y�$2"�!M��+ �@�@����X���iDU��0���
q���ϖ(��\���J�P/*�9 ��W�}��� ˘�-¨��,61f��n���`#E �G�PY�%�����a#�a��nx�2���
&Ȁ�&�A�f��F�1��N�D�0���7�`hǇ|�Y��lԔs������2�gi�$!=�d�C<!c�b�Q϶J��i�\\u�1
�Ԋ f��$1�bH��BX펒�:6g�U�W � �gi'P����*�Hd�5��C@�XB�\�_�AkaI^2JUA���?���x�`�2G�q��L30@�b�B4�6���-2�2.!��B�NW��rE8P��Nd