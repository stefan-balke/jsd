BZh91AY&SY	�Z� �߀Px���������P�oclv� P��U2M2� @4�h�h  J�T���~�oRi�2i�M0�2i�A�		4�5=OS�<Sj@��50�A�ޒh`LM&L�LM2100Q&�504�ɐ��i SC'��,�� DI�K)>=���ʗ� �B��XS_VmÍ�����aG��T����<�w>����,Ǉ!��S(��u�kۅ�נ\��P�r׋�����s};C�)8Q DG=��LĔ�QѦ�Ϊe^�5F��5�D!~8+P�����IR���K{o]K� `ǳ����ȍ�tN��Rmq�QN�[����f3Sb]�"|��}xҖj�K��鳑K��2B;e[�ãTl�+x���%k�
���B�>��B�Q(��jW��{5���cs�2��R�m��C�����R^S���
y�Q*Q%ʴ�ݜ\d��6�#rF�S�>�P�T(���
���Q�xL�P��R��]�.�_|�L2�"'9��9UU�仇��c�p`�0�c�ѷ{��zfKP�����U�X2�i$a* �9��Ơ��$#��R<
AC#K�{�1؊�ĩŕG�<�7�G�+�b#�ֺ#�<a��Q����l`u/6P��Β����q3ʒ|�
�3����à�����P��r�k�gpd[�B�����-f�o��Ϗ'2��	&�-��^]؟X�N����[3�-F��������n�q$�{�#�d9�����x��{u�][ag�o���fw�y�h��ϼ��a�^���0�B�#�a�9]uݜ7CZ����ɭ7��c�&뺓�2l���2Լ��rF�M3
Ջ��ɛr���X�h��F���(,A�Ą�h�B����_.	`��r������R��tZߓ���;o�=eD�����(z^U��}�84��S���.g��:٪��ja������|�Q0�%$���2-*��3/u=L����r��Ӳm�2�2�"�5���l0���qEԅg8�iq��
�V,���V���&h�lcBb�oZq��,/�'�m�jX��(e=�ol�5yN�M�(�Q��l3H�X���κUXX�Ƈ���o����W߼����@F�%�?x��)�Nr�x