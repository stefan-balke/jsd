BZh91AY&SY�h7 �_�Px����������P��;���4	�$�14bM2h2i��hd ���d� dh     HH���OS�SL#���a��M�0L@0	�h�h`ba"BhM2j�Oy="� ��y`�J 
�� ���~���A�DhT0$&S_ث�]�#a�dfX@>�EM�#���\y:=�9x�M:'u��g�
�V��q �R$D/l���|�*r+ L���rQy�YL'�6D���s<�{��3^P�-2��$jO!���9��%�� ֶ=Ol� V�bs�T�r���_�ͯ�O2�aHL32a��Ca
�8��)l
���Y.�u'Z�)XeK�;Y/J������Eaj���B�UZ�f��V�h%�h�2�f�%��Z��C[0�2W!JiJ��b"M8Jj�-�3��g���AOs Td5�mk�9��K�y��3A��V�@��`*�fɘ�HI�f(�7NF��~����0YY�D�V6�P�:3�	�]�'h(�,�H�	���b�2&�T�����&�Mp�8jUcw:�a���o�m��%t��;��P���9P��R�-��9UU%X�0�5�hǒ�*`�p�e6Sp�j����F]([TPP0�s�����7=�uT��4��DP�.p�5u���n���|�Svka��I��-%rg��^�LV�<x���Þ��������N	�A.��z���zC��C �#$/`r����Ƌ��*�tr�l��/!��ItJ��B���3<�I�07�j�L�n<�_��A��I<h��n�Bn�A���j*���wˋT@�q`����\�5�b����yY�C�>�'"ۥ%	��C���B����=.�6�)�e	��!�����P!uuP͌���#�Q��Y���3�5JhY���(�jk�&r_�טj����rB�R��@8�T~{���Zٯ~hh����6萼{΀4s)�?��:Ǥ5�#�
d�"s6������n (��PE�;�âB1�.�p�+��v����0��%,��i,�HME���P ŒQ'��.hC=��� ^�34=Ik8xL}a�hL���8�IW��@4<�V�`M�=��Y�Z�k�[�Pm;�3�D4H�ȄPx�e�8��F"�e����8�EI)v����(��/��!�����P;�U.��Am�A��%�2,@і�N摏�鉽��<H8u���4*f�,��h���ꦦ��h�Z���#��I�B���]��BC����