BZh91AY&SYE�V� �_�Py���������`z�աI�q* ������@�� ��  �220CFi�F i�# �������h @4� ��$�	=z�)�@  F��dd2`��&�F�@�&F I "i�LM&S��=LhMOD�����y�6/��4���L!�RE�W���UsH�N��b(1``�?���aJ��L����T��*�����j`�i�����ԫV��7NiũI$�n/��h�lv_�n�X�I��-'y�[�g���wzw�\��ӏ-w�d���ԫ��K:%M��_�M�c}��������s/T�����/H���DK6䉰9�kqL:��Y7/���*l
����}?�w�m��r�,����]s�9I��ʗ���dtn�Kȉu|\�-�c0��1��EI/2H吮��m���^d�Hc���ʩ,��/���gr�.iHf��Rȵ		iI|+A7�0�\���LX��)�2j�l����d��P��
3�K�M�1?f]p�־ƍ6�4�Gh��v*��L�^3��(�"�EU!�$�WT�lt��u��(�ٸ*�H$uy����*�LP��$vXj�,R:��I2H�J��u�R�Kd1��B�@BX�B0,`�����O~�r��>��Ɓ@�m���u������V1�;4 H�0�?~����|�����A�9~��EcU�<^�2��=DvXU�t�	�~D�>AūOv��ii>��q�A�H���y���7�笥�h{埶�O���<��9�yFOpS�&�p�UR��	�s��+��/��a�2�%��2�*�I�Wt ��뫒�-p(����-f$ޡ!H;ŻrΖ%�E�iE�6T��q0*SE�����[�K�e1��9��3F0�i�V��T��r�N������؟Z7�s��h��/K�Ք�������1X���J��}1��~�{Գ��1i6]���u�띌g#l���v������i�\p�r�l�"ŋo�>fK��Sڣn���M�uH:����=����c��U',Mo��McVIԼxiha�Y�Jk�����Sj�I%,�R��3|���,��{���Z�J���]l�f�f�k;JZ���2L"�5+3�f��R��)�9%u�!�z^	�v����G���6�~*?��^�,�\��n��s���G8��v�A�RO%�?�|�k�P[�7IQU�R���9����o����=�6��K���F���Xm Mz����D�~��D8�5��B��|�n�QL!	�,��aw�v`�VY����R�r���ۋF{3^g3R=.�3�/:2��+~=������Zt�}IP���W<WF�I�v���ke�Gs�g�~5R|��gFX�OΜ�x����1�!����)�,��