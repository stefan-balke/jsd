BZh91AY&SY��� S߀Px���������P^��.a��5ф�
��zLP��
�2���	� �F��~J��      HJhj���=56�@�z�  4�	���dɓ#	�i�F& �"@��%?I�T������=OP b4��S�^M y���Y���~㑨G�(X���e5�|p9��4,��0����PH�H|Z΍\��v�C���c�a��Nm?K�sw��D�aCno��;$8����-����i�b�����o�e�.7%>G�1.��5{Z�DHΙQ V����zG0�@�w�w��&�1�i�q�.苣1i��uA�T#��3馩V�G����TI64U�/�#Ir��|)����.�	r6���͙��x������E��cB(KDॕI��zbnP��UR��ZHV�v���*:�@+b*��"a9-fň<`���q�i�ʒR�ln5�lcwm��J����%�a�RNӒ�R�#��k#�L�F�#rF�`F�"q�b3-��da|T0����������)��r��<�W�)A�PH>��<2a�8��������x�<鷄e<�d�x풡�aVm?'z2������@ظ	��ш�.���ƥ�X`h��8�����3�2Ր���Aq��Խ&�\W�e�������D���,c�ʁaZ��6��(��fҁ��� �-�I<(�mu��'F���4�"�l��Ւe��&�0k�5�)XR�B��Ʒ���bƵ��@����� �73����`�Q��g>!��S�`b]�K��8U�M{췓 2�))�^�/Ē�-Q>dO@1_��B��M�Z`%U��/9�/�Z�\�g�0X���ݘ�wQ�G�#��eE�r�e�oEF�[s=AXnx�Q#�+� ��˱A(x�,HHF��H�\+u�X�T�!���T&��K=���	��!.��S���2zN��;���axHn�3���1;d?Xd4&W��8�$�,��8�o�L4�JG��YI�g*��VPFӒq�!���Hy��-y��0f��NN�~Ɍ^�j%�B�g�(]�C5��X���������$��\�%�ʠ����{ZE}�f�A���:3&%�L�گ,�"�@|s����-w���A���UX{���]��BB'߶@