BZh91AY&SYV0" �_�Py���������`�<@�9@� J!#M�=�~��A����z��4�4�J  �     8ɓ&# &L �# C ���7�   F�   2dɈ��	�����$H�53T��䧔�OQ�h�G���4���A$� P ~��r1H���B��I$�{� ��xMW�
ɖa	CRrQ��ռ����r}�N�{���l\��\9��ظs�����#��������7�L���r��KI���Rx�]f�t�G���>;�H�t �s�ay	�5IA���B��>�VOC昒Ak���%@���d!�c%
�0�R�H>8[��?�@������C%�B�M	���6R�TL9WPřє�tZ`CK�3��Nv�,R�x`�!S
3(J<Vf����ﲺ�2�l&�TP\W��2	��L�Z3��(�n����d�5qRbZƚ꒤��j���
���b!	(�2�*H,45uS�)͇6�K��Wt M�L)C�UhT)^SH,j��Ɛ��(���Xq���^������fK�W�pi���{`(N��hJ�dV+���x)T�����n�!l�L*u�[Q���yz�wci\^�4�8�m�o\n1�,�9���/UZ(�;]s=P޺���p�)���.Y&3�"�������ً.�"-L]��K"�*0��$EQ�
���ܲ�cr�#]3u�!KK@��LV���u2�n�ݢlQ8ln�/j)��4i7&�:Ј[�Q)�+������g�"^R�M'����ut��6Np����b#\6��Iv�P��ã�
���?��x��I�!�y���|D�H����h�F�	V�}���z
��RH<���Om��&o`m_�&��fØ�}�K ����$�J���DU\жz���6B(K��7�D&Q!s4s�g@��XE+
\�������υ������'9���������b�%1@P�q����Y&$��)��h�dt�/��P����YM7ݞҋhjS480�c�����箦�̒1Y�(���05k^��Pѥb�]w$���w �#%��l3�h96&E���X`P�jbS��+Ϛr�Dą�� $y�� �:J�!!��M�J�@�1�s�&H��*!"l`�hݐ���Oe"���o$H� 4�`��Y(dy% z9}r7�#"�Xl)��9�ĀE�yбB�0�ݵ$	�2g�J��Q�B��CHPm9�g$1�K$Lp��m��Fl�o�U�V�߀�F�H�:�ԝ�p(�
�H�3#J��ҁ����H-a�t��0E@d���J�cH��{uf�Iu�q�l��H��فQ,��7o���sk�nT���dn!#1�B�����H�
��@