BZh91AY&SYZ��� �_�Px���������`��ˊ�@��I MS�OJl�2x��h�?T�LCMhdѵ� �J?R'�Dh�4�&	�a � �`�2��j��*2!�i���#Ci�1 � �`�2��H�$Ѡ���I��6H� hi��ڌ�:!!�$�*�J�B����`��ci��d��=�m��a�Xf�9�'" h���e�����9�uz�n����9�ֵ/�b��趕����E���a��G<�:<b#��,$�r�֣��Er0`6�*���'�
:_ ~��|����Ðsu�1"���D�C�J����A���<f��Nlռ�%ܮ(���%����;$� �6�e��g ��ͭ9�cvԧ�	A��K{ԅB]�hT����	���ǯx@:/Y����ܭ�S�-�7��D�!8QƗe��
h��8�v�:�饘���N��g�p+�U�2�RUeTA�b4�����rg��q�6��-�a��*�R�S4�-)Sjn�+7�å��Z�[%٥�қ2�Fk[��Xrռ�W�:ᤫ@Q�$�6��T�դ�&-�轰j�с�p�XU<ʎ\p�|].>�U�5�3E�dX�\;�NB�.c�n+}
�į�>c����7�m���"7��>@�˛/�7bTS�����*̔�e	99�6�`�b i"g9 	  �h"6C�'�P	L�r5	���M��.�Le%|��JA aq�Ζ6L� ��Ռs��k�������}u�:9BA��'NN��л{?�P��q���@9���"xobhz�i��Rk�f�g7��,ǽ�ga���+z��nz�p���/���Pw{�@j�#<��¸�`=��n�+���c�OΒ��V� �Dc�I��2h,�y܊&!�J����E��bQ�mMI�4��67hPb�E	v߾AD�@F��֘!�L�)XT'T�q�l_�!�|�ʫ�ͦ�i�1�q��U�b"�������a��V�	��D=f��=�``�z/�C��$h�HM_����Te�FHY[���VdQAh&u/�������5�b:��m`@@G�4q��n{2���iZ�!Y팀G��� ���,z���A�R�jE*@�
� 	�jf���Q��HY�
̴JH(@�]1Ȉ!��	U"��%f3"��g��&����A6D���HOu>&�f��ILhy��OG���X8@�� ���N�tpb4&[��8��t����;A�\�� �a"i3�֯,z�9��z��i�7�$@1I�$:��wёQ�v�V�V������X�BjO5�� ����牀`�I�K�*�DxNc%����=IB�Gid�w5
�&�ȃ��=�s�S&b��E���#�(���	fUO�}�N6�A�`d,zw�e����"�(H-�� 