BZh91AY&SY(�' �߀Px���������`�
�<g@  %T���&C@ hɦ@  �	��2 ��@�   sbh0�2d��`�i���!�i�$��� M4�&�@ ���&L�20�&�db``$&@Ba�2z��h I��bM!�$  �V�HD����Y&�A�hR��@A&��pS+ƅ`e�BCGsR���+B�g��7�w�p���/.�����ҳ.��֗D�l�tq�L�;��OLU^�ޅ3K��r�d�;�"��C�N��sB�]����Ɨȡ�.37�8�`�fa�d慻(t��#%���0I���QVJ�_�6@�<P0����4���Ĥ���}��H`ǆ�`xw�����e�dc��vf8fs�0�p[��E
��R�^�)�N���%"��6��]��ơp�D�1��FԪ���F�"(BQ�D˲��� E�d�$@�ܑ F��U�C"I�ć�L:�U���C�«�)%����fr��1��#��E��
3`�L>T4�`U$:���
�F��ƛY4�M��l�Yʲ�xAh-�*�15������P��v`��.nl�e�x��kn��4#m���i&��DX�/b�<.ت|�2�d8�W�q� J!p ��I��וֹ�mLG%��-L(*we9r��M�*lT��j¶�Ù�b�V��\&�����%"�6����reNP��JA aaֶ�I�!��_�M����u{˭�����Pނ.(*���A|jRnz���&Na�x��Ve6��z���[9D�m� :w� ���LAms�I�z7�.�O�?�{��%}F$�B��q�^:�0��!v�����x��HV�_��Iy�AT�}bA�L�|�7�7/�J�L�l(g�� �-�I<��mvh��n慬��bY�62B]XG3TBef���:DL��U�)YG��5��z�+�!!�i0*���oP��X�����J��&P�#�?�t�H:$4�I��*��E}�v��[*��Jh[v���$ɞ� �>ys�4|��j��$�d��(м��#�Zח�h�g���:�������`�-���5i.%4��ɆLJs5a���D!M@:u( ��bdAC��d�(�@�%6oa�eI�* "&Ȁ�w�A�pB{)�H>��s����f ��|��`�37���q�>�ř�c�cBe}a�$��@G��G-�A�&�3�J���;K��Wu�4Ӛq�2C&1����X�h�ņm�͠U�W�֑b�
)���PH*c""�a��4BC�s�a��놅�RZ֠�����>M#?�ᙽ��^���`^�څ"�ՁQ-;��G7*b��-w��#A�`Я�;u�w$S�	��p