BZh91AY&SY�}�� �_�Px����������P�7N�eܩ���(�z�Se2�Ѡ2dS5�h4�@���(TzG��7�bh�I�10 i��JiCA��z�h�    *4 ~��  �   *H��h�6&B2j3F�� �a4��+��-c3�d+����w ��D���"���?�*�Ƿ53�£�R�Z�&v���:�\0��L{O�T���Wm~�l+Z�@�Ο���sT�O�aGu�5H�o%��	}��ϺU�Ш�E��4���28<�)�$飱�E���qo�pZ��f�|L��Aq�����!�rӱU�#�����0����$���2(bX��n�7L�\��5��Q%�EkL��-xh�9�c�f�������յi��S�逄�(P��]�;��♾�Ưbe�X�y���.��,K���oES���r�*�'X(֕��C��༲kM�����}Xt5��ga�p�F��L�-0L�úW�w&ٶ�Ԕ�� �V���m@���~��v1���t�8Z��ERR���OV��k�4��$!,��I@� c0T\�Io�9d�
��\��EA"P�B%�᫈��
�%�AN�T�2���
�o���a{.,�+�\��:f���DU���*��e���trɊs	��hh��L��a��M�^�p���%Е��_5y5#Q�\讱gu0����;�xy(�N.����$z·O>4ǜ?�98�!����b^s50�F��-�|���l�ς�v�L{�IRG�����Js��=יĥ�����z)c��c3.V��~�F��;�˦s��a�kZ�R E�,���Zt���>4�e�*�{��f��UEI*�غy�̼��EnѰ�8�5�R�K������^�H��Ų��v��c��?���u�q��K�mqմ5/�i8������}�ѱt�D/܂R��*�x��Y<瞮}�I�5ci��#��G��j�z����f.Vk�FJ�J&5�Z�XV��kt�D�+^E���;�f,	�t��S��&)z���b[
ZŴ��:�D�l|)�NW"T���3���9"ã�͍��57�ث��TJg��ג+�kEGJ9�R5�H���43u��#�8�y9�R��8pR�Ty���h�X��H׾����>T�їÌip���da/Z8��Q���8bgd�|�U����"THԩV" �H�6����z��J\o�l4T6Ȼ6��Ț�o�u�^�5Sڼ�s��I�@�PTH�rE8P��}��