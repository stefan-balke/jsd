BZh91AY&SYe�Y �_�Px����������`}w�O]	A��|{@h5P�M6���z�C�2A�A�M��)4 �   2   ��MT��=F�M �   @!!!��=@�   h �T�O���F�ځ��   h *I	�`�I�$�����4 �2i��|��2HZD�K!^�w櫖��YD��5|�h��F8�2�c)��*9T��D1�ˌ��������q��.z�D�L��g\L#b5�����Q�\*�E�D�BvK	)�ٿH���̯|`�,�(�Y�$�X��� �7�<�X�̍&��lיi�#��2Mocr�$%%ʀ�К��㾲�A �mw�T \	#�@)J����a��;*�ͻ`�B�8��\�ƓO3K��KKm�,�<�Y	����{K�e��
Q���6tk�(�:�a �y�O����5�FU����Ŕi}5�y) L�<H\!`P�7����g&[�kI�0ȗ��cHu$"h�n�S���YA�^��&\/P���r�����+���4�ʬ0}p�s�BMY/,�.�D�X�� � B����K�*�1(�����t�BQ�.�di�T%���)����	ژ���EY1lY�v�.Q���04@z�L.�<,0�Ȃ­M2�cYQt���+�Iʍ9"-%�0�7fcN�d���+d@��d6�X%�.�WT�B/aw3%�W�7� �A��m$�C��th\|$r�I!�qQ*Q%�b�)�P���1����ccc�4l���A2��$nʪ�Q8B1�B�2�V�hb�
��>|���W#Λ����F8�W#e��x�w�B��p�	�y�N�g3��́�F��8��:!m���w�%����UT�7�}�֦�_s�#���*FE���$��<Oc��L�zυ�g�L۔�?�б�gy���nѵ08�,?���$_��{���I�G�d��'zH�j�׿S}��t�%-M��C����=��i%j��&L���)H�X
�M���mP*$�S RXà�Hen��R���O+:X���L��O�"�*��9:��L~uz���sn:\�����O���a��r�$���Q|�]c��'�۱ҽr�#r-/�&��y�_;�L�-[���9����9�M�%��^��hW>L�4p�4�XZD�Gg��Tu�񫺮��3�ib�JF
W��,%�oQ�m�Ȥ$�n�PE˔9��D�`/a!t�����1�Y[�ꌇ��K_KX�}�����aВ;\H�SKA%�����q=:[f����k|�F蚝=�+�ب�ǭ�u��Ex�"���M�#Y|�{�fb�x�N����f�dUJ���K��*��Z/V�M\-ł�w�Ҝ��s����-�1/�V}LFF{�������hT�]S�!Ց����^nP�
���b����W�R���>��\[L��E�[�3 ���6
t��t語�	�;�y�zt*�TL����w$S�	 &]�