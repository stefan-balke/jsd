BZh91AY&SY
�� �߀Px����������P�wYmQ�  Ji��ڃC�d�&��`2�E ѣM ���h %=D��MM�Q�����a=F� �hs F	�0M`�L$H $�hMOS���P=@4S�a��I>��	"�j@������h@}!Z� ���5�?ɸ" <�."�]	!���h�"̆G����fկ?j��'q��Fe_a�@�4r.]ϔ�������MP��s>+U�����ڽ�d��acG�w{�͘cl�������}ċӸ��j�)�)L��6T�����Z��|� ���!!P+�b�ŭ0�3�K���o�b�d��995�;���~�ڡt�HM
o�R0��� �L2�`�����Kg�/*�ġ��ҚR�
�7(f��SPL���mJ@�"�g4m��ߙ�a�ɕŐ/!�"��[ШX�z������) V4/�x�J��	�3�CR�m���!p�0F��1�Z��&�J���(D�L:�P�gn����H;#j	��Ѝ�z:�#..��M"��.eU`b�N>�<�G/��q��
�.b�R�$UT㵋3=U4"��QIH"6&Q��	a-R(�-��
%�SJB�@�ez��K��>|1�_6���,>�����@ 5�e�c����!�W ��!H��-�77��t`�SL��n��ց�Ȗ�Qbb�;�z�W�����i��� ��}�xf)�h2h�/~3�_1�nIzt����0l>�
��`k_+&��fe��� �,����)J�-�,�h39������El)�� eX�q&�3�D��{�y	E�LlMW�@ȝX6�"p�£
�98��Ӡ� {��-Eƕ1@P�����k�R`�.Y�K�IuGG���n��yBF��YMc�׸��
f�0e��5��f��3�n�f�@@G"��Mk^��Pѡp4�g]�Y�G%z��K:
�4�
�"s2
�s���hy @H��@��+1Ȉ!��"
$A@�"��2��ʓD4T> �M��܅��By�P��p�`3Aۈ��d��G��x}�M�A c���o;����XЙNc��[�i4�����``×�p��&���yi�t����P�(6��3��� ң�Hw��lo(3=��a�7�-�$XN�5'u�E*�Ȉn �b��Ӥ�pԺ����9IpB�T�>r���^�cI�xs{Ak4,3W�H�v�-�6�3j����d4��+1=�W�rE8P�
��