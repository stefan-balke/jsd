BZh91AY&SY��� '߀Px���������P�!#0ѓ@Q)��4��)�=@� =@  h9�14L�2da0M4����$B T�@�=O(� @ �h`LM&L�LM2100	4��M2���5<��@4d�SB�Z! VHD6����hR�d��М89�B�hX��&�B�m �@\���ܹ��cW���d��p^Y$r�y,�=��'���;E�1�P�q2y�������T�1����<�3M=��� �>��Z�`�w�M +Y�H@��a�ZZe�O/�Z>e�L����E�-����f�q$�ݪ�4✩�\�p���pa���,針�C����G�x�X�m�FLM(�Ɏ�^LiB�9Dc��2��l�C%5$J���Q��t���D���K��"��l�"�F��k��L'{.�X�Eh�R�p���7���hhPA��m��R��!��"v��1$EZ��tܺ,���ķ&(mTCe��MBG(eLR��$��av�f�&4��i�WGC0l�ce�k�6��0����ҳ�`��5o�����O��<'�b�{��J*�1�þ�[UV�$�b��i����~&�����jWt�!!y��W���3H�{^-\��e���{�Dy�F,��
	���j�L�j*g{ ��[�I�J��L�F�1i:4�j�!'�8�Մ��lM f�g�*�Ո�g%l�=9���N1(}Z��^���ˮ5���A@l(X�a���M:S|�Y%��9�}�<����&@j��z�>�4���;%�G��� �L䂢0�4@'�$��t�T��>KAyv�4r�Sa����s�%�ň���9�B���NQ�4�� @H�ҠD���D4��Y"��M����.M�P��� "�<W~�'����]F�@��gH��=��<�l0��#��Y�Ph)�t��Đ��3	�����8�b�\UŎ������P�(6��3v��%X�&8�Xl��Fkٷ0��P�*�m���:�)���(
�Y�i0XP�a@���H�-��&A����¢���4���fc���� ��4��b�cR�U,u�D��p:^��-��f&�k4,��˩���"�(H	L�X 