BZh91AY&SYk�`� (߀Px����������P>s�v��	 p�H�=#�=T�=OSM24�h�C  hhh%LCD���@ h�  h �ȉ5O�4��4Ї��hѠs F	�0M`�L$HхI��=O�Q� @�M=&�`���IPH,!@����1ȽAV�$�&�d�����p/9�+��d�0b�Z�R7 `�b�����Ɔ��ޮ���oM�dJ$}ϭ�R5^1]�B�uJP��S�Ϝ�J�G�j]�%����Ą&RD��ʊY�Z1���eJm�OU;Pb�����m�U�O���|��F<�,	&L4��0;�U�č�٢�B�e��~sC���tCFWE��U4��6/&��/MaD:�Qn���g:��y:���󳽃��"֓R�Jq ����L���M	��]�@�F�QY�JR-�r�*��3�^D�Ua��aQ�F|:Μ�ڵx6�B�I$�� 1�tv���#f���Q%��N��^��UXU�NK�Z��Pچ���Ш��¢�,1�V2HH j4䍱A	BA�1��D��\T�Gɳk,�È$�[���F��ۜe��(Y�KA3<^�a��*�Kr^.ʢ}n�\ �
J�°��f
�b��/pr�Jp�#,,�'��0�B�(G�H�);���Tx���dͧ�@�L��ؽ�Jl�C6��}^�3GrI�@�ku�2zk:��Р��DP�\Z�2�3L��K�!�Zb��*��Κ�C���E���i��m�:5�����{��ƃ%1@P�g0b�|�̜��u�b5�D�R#~��0�$C�=&D�F��T��=dn�e�SP�����R\n�mh�pֽ7��V�ǆ�1`��\�^]�x%:�����q��P``L/h�̂��񛼐��@:2L�B���P�ljx�X1!X#t���5;�,%�6D_���ބ�SZK��0�zG�ŞV��:>x6�~'���k+�x�� >�1� �f�A0�钸���4h��.�*6�3<�Hcte(DǬ�o�ʌۻ<EXEt�zr3���MIݧ�D�M2nA�//CP)5�P�SE�$����%�U@�FQ���cH����mi1yg��.h6��V���H������י�R����!�k4+-)�.�p� ����