BZh91AY&SY�D �_�Py���������P�.�V�`
 	DA��	=4��zA�z�h4  &LBS@ d     	L��@� 4    ��2b10d�2 h�00I#Bd�@ML	=M�M!�@l�yM���;�%��e�|夌H�����	J��Z&UU$�T��f
4|oUV,`jTQ�Rz�aURFv����*��my�]��)�v^�H 5��4g�S��T��E��P%4!%8�rJ������xwt�&�e)���X��l�%Ru��G��f�|}q7�5���$I��V8�L�G��׾O�橅�9Uf��q�Թ�*RR�����u�Th�6�tb3g�����%$<�h�N��{�P����J���i�F��ەI-G�E�W-mR�F�`j�P�#zSX0���H��	���3RII(
�\F�J�겖2���%�A����H���3{+��p���,
l��JL��34L�������"൳�Lڴb�Ok�T�R�[�UUUE@�_�/l��LA�i%��w�r��ʄ�V	D��m"�D|MB�L���X����(���P�%���rL�T�Q�
���G�cj��vftc��+����S�=�����$qjP`&�')݌q�ڴH�/k���*�т�łq�kKJ�2 L�gxi�a!���Û�z���=P�ʠ��i7���[8�'4����Y:.>3�mf�O�TӲ��(����~�K���S��g$�����꥖|��V�e��.�V�8��6T��Y�KE�x���S\R��N�BS�F%�_+L2[ڧ�-�U��S6��*IVt.��32�+w��W#�I�p.�0z������)(<0X�g&�`��G�œ�M?6���%��%Fxc$���>�����aP*E�%t����y
@*�D��bŶϟ#b�d�'��9�Rn��I;��`}��z�Q���S�Tr\�؝��;%{�����3�V<1an�2�B���X�LK�VY����T>^%�iv9T�)���ɌYQ��d���م�nv�O��$�w��I�)���S�����>�s{��,OG���͹~�y�
�S���Σ6W|��Rx�)<=\à�b��ML�3��xCG�I���V0��ڦ
S��LUmgR��k;��ϳjd�e����S�<�.̼Ƶ��\2pon^b����7��-k��i�E0��P�c���U�G
����'��u�tԔ��a<�.��D�0hэ5��Y��c��Ҩ�:���N�H�QRJ�O�]��B@S��