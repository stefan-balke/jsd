BZh91AY&SY� �_�Px���������P��NZT���$�5A�M=@�F��hi�����S@Q�� �B$�5M�O5Ci<���S� ���A�ɓ&F�L�LRHa2bb���=O&���  4��4/�+��-a2�d+��}깦�(��D���X��k���p=v7)3, 4z�JF́����w���R0Z�𬘱�# �ݑ�Ki���+�o�|��L����X�����>^@���6h3&��	��5O��c����!��:dq:��֝��BI��$+!&��S�h�{O�R�*Q�MѪ;�ǆ!!���\�F��m�^��r����63w0h8��St��z�*���P�@�����3��v����J �(L�k{����S4���Ix7g5
�S�L-��jP�B-)ْQX�(�$�M�Y����`I�V��8�P��3Y��Î�^�'��Q�a�6l�z�2\P���]��9�jB�,�l۫�cVE�upnRP�Y@��c�_�	a$���D!��}�夻��B�'��R�/y �YM\��FrB�L���,ES�H��]@�AօA@�5ڶ�@�l[x=�������k���yC���xǞ}:�.՘p�k�Y����Q!�$�=#�&�����#�.>A�咖��ff��#Z��G��0�Z�h��h0P�0�ځ�p[	��)��F�@qQ�N�y}�e�I��4���H�/F˛���;�]-R_=��a����K,��w�5�����u݁x��H�>���P�dF
��=ְ��$rM#��C�E�[�4������!ٯ2��{�l�Nu�DU�']��E���5�ǚ�I���蘥�K�����ٲQI��O�tj�=_=�m���q��.�&��w���o0��������o4���vjnH�g�7Q,X���n4+f=��������k��ʬx�sw;�G[�zꍸޓ^�K��*��L.�p�7�7S�hA��(�s�"��<i,����YXH��+Fr�ݱ_���b%���[GN�ÄJۇBG�ȼSS٨.R<��{r>}M�%�W��#{��J���+�mTJa��r2]$WP�EG�YG_w���0Y��d���z�^�x`m;@��eg�%"�0am&��3)�����ю��sK�W2_�|����0HŞ�-k6��&�K&�Zpdr�3�θ3��v��a/�_KH��>\�SI�����jd\ɶgbMwE�8��xh���L��ib� ���-��.�p� 866