BZh91AY&SY��@T p_�Px����������P�r$���� R�&�e='꟤���h�I�� 444�MiQ� Ѡ F@  �H�����4�ɦ�O)�hLЁ�#@i��� �`�2��H� L���I���zOP@6����M|�	$��$(>���9 <!Z���$���fہw�I^4+&\���Ңdhn.l,�`g���͹�f�ÿ罚�[��H������(��` i�$��6A+Q/	A��>Cs1��bf����F)�8�b=	��+9��d�x=�HB��_J!
�r_�6&8��o	ȭ�{��#��˨��Bɗ��!����Z�l���5�FZ+�]p�R$Ja5,;�؄HK�[_�+����諴�0z�ХtM���rsUhsT�|��)0�jIR�u�s�b�جMBl�UeF�٢xʪ���J�,Y(]l��(X�Af+�j�QTR���$��B�ADUq���hPK���JtyY��9�$P����J 1�T6t�䑫HӖH
��G.F�(�~�c�Q�Z��%$*@�r�n)1�$QIai����	k���L�^�9'��Ǻ�����F��yK�y�k��!/��&�:{�Hh�!e�1ω���W2������fJQ'N;��GKE�3Fa�5J�Z����Ă�������G��[E@�,H�	��_L@����),hhьIs iD�}�� ��䉌j��}�l���ZI�@�ku�؇sq�ۋvj�E�%Ū �ȘZ!��@�FG\�:Eq�x�f{t8���Xֱ� Ƅ�iC��X+��w�=��g �`kTIu�����T�������Mz	#n4o�k��L�SP�|hb%�$'����F�Bu5�3���>��m��7�q�%���pj���]k\�7�ũgHB[8 wz��<�:��r��@��feĹR��̘jh'2�Xny��I$� 	�( ���94�$Q"�xNl�Z�5:��*���"1�=���l �9�0��
��e��iG+�
�,����~�AMm�6F!2��yĐ�5�р1�2=< 4
3�Eyc��C�����FӢq�H�iz�i���f��Ĩ���sa�8��6�bu	�;��(S	����1�K#.b���o$���n���J�b�F��^�����hoi1�n�p^�oE���3� ���r��;�EKZ�{4���E����)�<�