BZh91AY&SY�_> _�Px���������P�֩E$����h�d�h��CF��A�ɓ&F�L�LBAMHi�F�������  i�`LM&L�LM2100	�Ƃ	��H���44 �z&��i'�!�� ! ~?�r4�,5$XC)�q}�ۇ5�Z#2�&�6���2i8wM}���|���32չL�sm�.��oG��-�;J��/Ҷ�N��Z�!��mfy�Q�/5n��H�5�(=$��;���X�=\i�h�$K,�H h-�ZH.��4y��*�_�@���c㟿�9{!���9imZU"��QNR��F�2�����_c-%�gXɃ�U��DbE�
�}p�F#U�vR��\��4!P�jfK�lձ.����rErj��+s������TB��KI��-��WY콥&����0���lccѶ�hi�'p���K��G*�y�D�D��K��ԵSd��~eg������H�e�FaBڨ��a��]F6&����:�������.��;u�,wr����=F��v�Sfy�9M�(�*���<,�	��5]��X��f�fuʗ�VR[��rGpU����(~�0c�F�r����;!D�
 �9��L��V���I-�I�#"q��N)?#	���|�B�!���r�dx�Ғz��n��F���`U�6�B]w���Q�X�&a�)T��t�8��4��`C@�"��`��~�5�~�s)���N���)�I�� �3��k��:#��v]n�odj��Jh[_v���f�C�P�c��Ӹ4�˶��f"�kbn�a���j�y��z5,�����Dq��:J����@��2�X��T`j&X�3�+�)�5@���A���$$#��]"�xݛ�5���Dh�xL�c���:��B{��#�t��̏fB,L�I�w�vG�h	��>	�2<$>��4&W���BĒR�:����&��Y+̚f���:�`m:@��҈�����Z7F��6gv�V\~I��,N�5��a��,c""���4@��k,la��놎���J�����*��E��-&�KQ��<�Ʌ���cgP�K\��p�;2�/������ �02��r��.�p�!��|