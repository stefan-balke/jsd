BZh91AY&SYp6�� x߀Py����������`�y�ё 9������SFA� ��h   4)5@h4�z��2��8ɓM0�14`� Ѧ &��hPi�A�=A��@����4�	��0#F�` @�$h��	��5O5Oԙ�M��@Ѡ�є�֫�z$�2��!d+���́��F�IIX�M���n@fXD�G��RQ�  � b���7���]�ue�n�����Wv�p�UӺuwM.���;���;�د� ��(`|������E���������\�LH��J��M���KM�6���tw��u���vl�̚��|�m�j�"q�q �a��B����}6$�h�ժ� ���H�Nɣ�U����L��	URI$!8�[�����o����x� �>\���+.�\�����i�ͦc�B��uWU}��*:�ԃ�ɘ���Ҋr��c����H�����V�DI���҄N��Ȃk�\b4F���������WQ�Z�H�a�L)�wPk�F��pe��Azų���K���Q�\뗀3p���Ca��S[��;M�WZoU\)@	kr,�iw!ʒ z�3��!G	�˸U	�-�r]!�h�N��ס4�E���vHE'���YVn-4�f�$4d5�ކgJar��=�w�K�v3`�VW�z(rR�a��0�� ����x.B�d�� �b�s2�n]���5�n*X�Yv��r_r�Â�-UUH�q��*���(̚�z�X�9Jܶ�vVe�aa���k܎	��w��t�qOF��	�,��1^��ޢ�e�%��d���9f gLG4�Pl��^�p�Plcc��m�4�!��������B�C��T�KYj4��v+-��uC��,�]�HEm6w��M��i�ȍ������&	L)�����^&PՕu$�y�PP0�u>v��m$&ѳ�S��>�t��{�B��0H_?�K�Ap���I����A�Dv�8DA-�u��^YiQH���Rd��Ue�7�וI��w�'��):��'�=.�~S˵�?L=瘚x�������_cώ�	�2;�a�5�}rE�~��S�I&>�P�r/�7S�㑔��C����2�Z��ϖg��K,�4�I+m�2�N��R��4T��������y0��ՇJ�I�����LI2��0ki�"�z
��vgd83��8�ݰm6��Ns�`Z�~�Xg��6۫[znin�K0������7c�d��~NT�3ńt�=~��GlN���1�¿f�Nl�i�R����)�������������N��V+|�p:��,��ˌoY6M���B��@�~��*3_�^��˚�������t�5����	{���~5��� ��({}*����!�[�)Y���6�*��c��FG�̂���-��|�ϤJ�~��I��[Y%�#����h����&���=_f\]��NQ79꺼N
�L��n�l$��HޑQZ�l}]�d�B������tj4���9��\�U+(S�r�)ROe[oS"��Cgu�.�ޛ+FZN���]3����=���C}7!��p���� ͌�y��Z�T�몾�hی�8X���-��L|�F�r��*ܳ���i�q�0f�52fgw��S���;�zmT;TMZ����)����@