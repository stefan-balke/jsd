BZh91AY&SYC��� O߀Px���������P�wYXaÆڍ hJ$�&��4424i��4&�E4 4     �����z��4�OQ��  @4�	���dɓ#	�i�F& �"@��&Lf�ښ�mF�OQ�<�BhC� P�J�"��$����#��P�Uc��&���6��bJ�Y&HH�����R�L�ww����^���qyۧ�,G��#�O|�#��c��0Y��A�Z/wO9i������Væ������i5��F	�3��Р��9Ꙇ{��fZ^W͍����� V�y�Q+�2d����7��Uu�1XEݲ���t����
��{�	,��
}f���5^�+z���i�JI�Nv�M��8j��&�tF�>'-�@b�(RA*E ����fI^��*�R��55JN�2��Z`�ox��@��*L��R�R �)���V&�AX�!�A$��,�_lc�lEt*� 2'p��Jކ׺.E^-a��9��b�6.SM���+�a�ű#V�PI,�$̙T�0���G"`L!�D��TKxS�����iS�Q�9�{�_�D��a��PFwbCM=����P�|RFu�-܀3h�x�6G(O(U�i�~�H�aI]r��X� ŗ�q�p�υ��x�`��0]ݶ���<Bq"�����$0�B�(������A�1F���m�/<C��!y�N���t�,Љ0WW�FcP�EC����M�DR��j�c�N�ը52B]W�Q��t����%[B��6�ۑ��	�?[��#�;l0���3Ќ�R�HCpnP&�����'F����N�ǩ�t�$j	.�H�Tq��.հ��]��{\�T���9+Bdi|^���)'�Յ��4ܔ��85��:M���G�֯-h�pB4-0	\������GQ�,el5�Px-��b���2�X�5��s�9E��J�#$��sf��
�
���D�)�UR �0	ٛF\s;n(�4X/, �l�q�kv�۵	뮠{N���0�E�Αy2tz�z��>7.F!!�{�ty��N�}��hL���=Ab[�N�)�!^[ 3��3�ΰ,v�w�#�^v2��*6H�y"�p�a�f���K�k�Z\nSm�X�Ba��a�qP$�I�g-f`�F,���,-�J�� ���%,��H4|
�4��<�;I����8�)@��P�F�5K��B$�B�/05�5T�:�|7�Ӷa��4,x�=�+���"�(H!��� 