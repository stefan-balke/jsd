BZh91AY&SY+��? �_�Px����������P�r.�35F�4)=�16��S@��=G���C� �yA������       )�$jdjzO)�2i����    9�#� �&���0F&$Љ���&z���)� ��E(҄($ �B+I(�w`�2���Z��"k�_�py�@b4,���*6���AFF���k�pjע�~9��%�s��<�3�̈́Dߋ�z؍�V*e�F��!�'�r3z�
���~�����EK�bf�ұ|H.��T��2'	m���ރ%���b�g��U��1{�c���4�OT��˴�=oB���f�m���۳^�n��q�qҗ�K��@��H�m�I(4��k���t�"�C�Je ����ŨsL�c�����{��.3�Z3�],��z��b�	�Z�Ѡ9��+{�@u�(���k �@�b����Pqt+�"���ْ�!�K�Q�abs$\�U
̕,2�|t��X12Σ�
��Xj�W*�39�]�9�lcc��m�*(c:,uv��V�N2U+��8�ݯwR�~#�LX*�^B���$��Dq"6��9��V�1��e��,�sI��M�������ʹ�+�&��B����?��?qA^�g�e���a��\V����ʕ[#����m�6� ��N�\�Us�g0B:I�ǭk����Y�0G� �hH�q�L�DT �A y�9%=ޥ���K�YY4�z��Zɟ؄Rf�uh)ccPd�����A��1�I=u	Z�ކ��in;v�j�E�˓TI�H�c�]5x�aJ�<Y�\��g�YcE�x�Chhk(�0
­C�A��LW�,H�����{o�;'�@0GWU��Hd.�H�;{+��[↉QJ�>B+@fT�JO 3'�	w�)�����}K�������Ţ�H@8<�ϐ������6�1=A�b8��Ba�s5�a��̒@]@:5�Q��XPlhQ	z��K#I���ju()4T=����"2�|���lv��f�`�i����ۡ�f���ƻև�c��BezOY�,I} jE��:���a4�P���L���:E�UC�D�^����=�aqhoQq:uh*�+�r��r���MA(���A/!�C7��F��ԅ=jK�C ��e��.��FK�U h��M#1o�㉤�b@���ґcz�P5�q���ɵ�pT�����h6�/f���)�_�1�