BZh91AY&SY_8n  �߀Px����������P�����lq�Re�G	D&MOI��OML��Q�M�̧���@@�M$�@@    � ��e2I�� �4 h�& �4d40	�10�!4�4О�{T����Ꞡ�F�1ѨښI�1� PT^�$H@�>��I���B�i+ M}���ŒK1�`�4xZ���7��6uwz�9z�����Ц��
cSTh������Ҁ�5ɍ�c�Tb���~-��:8VeFT��s�4� �</ ՁJ���gD�^�9�!WF,�� P�fX�Я��e �F(�d�ENx����:�A2�
�
.L��yCz��l��"^���J.r�h6J
�+�DSCbv,4�$bn!'�0Z���3��j�7-W2����UXVXň��Pd[��9њ��ףՋ��M	�aEi7��Q!�M���5��K�aV�Uw6�&`�jp���K��	@�\*���N&Լ�԰1i��nQE1z�R�2���v�L��61��m�� �雼ᲅ��#�
�7��(���:���F�9j�m\dȄġӑ�)�]�PՊ��(Z��(F���A���h���&��z��¼��l��Vr�}l��#F��E��q0����	T�M+�0���R�c�j��*�c9�1`&��ΐ&Z z�&�ޚ����j�a�?��I���^Z����*T�5�6�
�=��X�%�3vi+�j������3(�V$����jD��|�WFA�o�pģU���kMZ���ը6�9�,ڠ���A�IA.��)������G{8�[�C><�K�ވ�l(�� �/ ,�z�`�I4x��u���c<T@r�C{�
.�h���:���M�x �V�L�I���&�M�AI��*���Qz�Ir�0�����!se!W�䘯XR�;������N��r�ʋ�s�E�a{A9�!��7����@�o9A �ŇD�h=��# �*���v��̅M1��Y�ږ��wpByt+���T��@�<��MC�e�R�^`IY���&*��7�RB�������:�;� ���h*s;C��NV�A`�t@��!���D��Ea�W���e�=b�e���I�(�k��<��d���p�H�7X�5�P3�WEIj09�M��d�P4`���CH���y���T}䎮fй��	2�4� �H��P���ꕭ��:A�`д��.�p� �p�@