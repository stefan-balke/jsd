BZh91AY&SY[5
 �_�Px���������`��^�Z\�  �xI�F�  hѦ�   5<�4JL���     9�14L�2da0M4����%=H���  4     �A�ɓ&F�L�LDBM4dhL���	� �A�2d���>"@@�J���_��?���95�_(Af� Њ!%��?�6�<h�+ƅrsHh�jd!���t@^�:Cw#Ow�T���{��%s�m��m�m�C�J%�GÏ����;-]�TŔʒ1�'��:|E��eA6�vI��?�q����sHִ�A8GG��	5'���I����)���
S�F+k��D���t�Z�J���m�Ӆ�^on�R�D9]�����!i�V�wX{<!�p�-��梵9��GRnt�j���V�S��������N��k>���6T���"G���"e����o	��q5������J!2(H����kX�+vK)(ॐ/�Á�� ;���.���C�%_*:�
q��8�^`f-��C#'*�$8V��w���;Z���c��E�Z��s�u�!shѧ�zV�58$MCZFC��f`4� �Q	� �*
'��`d:��P����P�S,���]���#CO;Tv�����`��'!E�-Kf˘��p�(����	I����锼:�q0H��y䉉")Z:� ��bf�%)2��JĲ���̋��J!x�P�
*�R��A*L�
_*BA�5ְ�B l��t�����14����#! o�ã�}���!ҭ��,{<)�x%��&B���� �l��85s0�S�&�k����
����<����~�I_�4 ��@d��g�b�oBr���	gԾ#.����M���A�FL�|�T����|nH�c!����dx�<�'�Bmm���k3;6�oCPnd"��aZ��*����&�3�E�1[B�)r���7jC����r�@8�Uto�؏�|��nh2TI������`Ѓ�C2WA(�du����!gd4Vh����yU�5�c�T�0�c��5����oB}:������G��|P��u��qCF+& [��1�<�4t���l3�i:�,K��a��@��T���Kuʓ(X(N��HP���B �!��"*�P�&��2�҅�",Yd�E��$�d'�v�i� f�ӭ ���O���n'X@�>�7q�zPJ[�3-�v@�� |�b	��������[
�=�A�v���u�5�FӢr�I �U�$q�Kh�Xf�u
Ћi:Pk8�%�,R��ȪX�#pC6����jp*j��A!u��+:��� (_-��*w4����#�I�{H:���{x����%�YJ*Iǔ�+�_��V����Ȅ��N�����"�(H-�� 