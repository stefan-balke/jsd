BZh91AY&SY�
b@ �߀Px���������P��՝Up�FB���O
O����Ї��d� �22dOI�"�  �   !!	� i�jd 4    sbh0�2d��`�i���!�*I h��MOA6�'�  �����-"�F2Id+���*�j�_��
���!����ٷ����hYɄ���Q#IH>=�������o��cћvj���'�{�pݺah��E���\�Z��ʮۅ�`R�+�m�WI��+�)����WP���"�H��I���kM�Z�k+]�c�U}�c����r�VU�Ï���Ȇ�!�M�;��S�J��^�OS�Fyu-T��(�!N���iX���7`���V�[�<,)�1���(��F4P-���ld0@Ij2�\��P
��̈EZ�q!�3S*x���1N��kIY;P8H��b1�9�4�+R)&�jֆY�-Ar�(�<�(_<�u������o��Z�nM�!�ؽK�[	ԭ�^.Z�V��r���������m��CB!�X��v���#�
�;tJ�Ik��h�e�mϾ-D�dk7���:M�۔866��e�4���PP0�q�w��&aU�j�����tKQFŕg�Ѭ �O	��<|���ŏ$��v��fЮyO>���#���^���>�A�S78M��78MM�P�t�L�hZ7��߁ꑟ�D��ca��]�ڷ%�iKNɹdۘ��$a�1�xj	�#�6����fJrP�>LbR���w}4��{L���]���aEg�nu�51�f�Z3.��Z��\�8B�"���|EX'��L5EYO���)��Ym�΍�&�����S�&PZ�'G�8���6ژ��x�������ZB���/�3D�#$,M��+d��^�)��gO!���Ë'5��"ŋj��*ۆz9x�\ʠnÐ�o3�*:Xu��7�4�����F
�ʤ_s�1�6�9��R�r�(,A�Ą�i�]"�V�3!��"4`=�-}(�M�����n#��/�͏f�%�G����v�#"���g�������nTL�1�u��+�lEGQJ2�q��^��SC��v4Iׁ�z�V�3��ee�yH����i����E��l9����~��ѧ���n�YM�sY�R��f9�1ѝq�*G[5�6ʹ�(�]��MH��\�u%�g���h��1p�XH�tY��c��UT�9&ls�T��ZTM9L�ܑN$%� 