BZh91AY&SY9x�� �߀Px���������P�ws7fA��P��S�i�=ODhd� h2=#�4hA��A�    h %2$Д�ODѦ4�14z�  �`LM&L�LM2100I@��2jMQ��=@CC i�Ml!+�D��c"3�K!_���*�{��%���{S�ª���A�RL�^ Ps(����K��k���ŷ¸�8>3|��˻R�Z��;�I��3H1��*��0����db�nT��$���W\hL1T�P0�#�B��hw(�R���/��`���@c��M��#ֶ��X@��^�aӱ��g����T�o�v����bc2�UWwd�8Fo�/��a(*
.!"j�D|�֦MR�nV��y1���nd�� �1£=-�,�e��+ǙH�n�J3�L2�3&�!"�. ��k�R�J"�©J2a7\�q!��dE(�`�[LV&&�upEC�j e(�y���׺�&�"E��T�g�t�-�����%�$�P( c9��tLF�cNY$
ϞG.F�ָ��
P鹧3GS�K���]��L�B&�!K�9B�*�HH j8�F��#>��R���N8l1���w~�pW�c.x��0��dڪtRr[>p��47O��E�r����QSSJ���z@4���G}g.�>3��?�}��F�����Ʒ�^n�})��R��q�φ�p�M��!�1�:)��bb��C�{o3�KS���/�j�8a|t�1d�L��]�7��5[��(�.��RE;��SU����-�N���YOo�6٧�%�Q*�ػx�x�������hd�1K�/�|����|���\��׎̣ÿ/�h�ɂ�GJі��^\z��ك����S_�woY���ǧs��;'�bŵ�+�cR��3�?|��l�P8ȅO���e�+}Q�S�f߹��$f�����a����Xo����A�ab�WD�.(b���ƢX�X2	��.*�j��6IW^���%p��#�v6���%ԏ��3>�������g�*6����:U�w<�k�Wh�
��l�z��`���K7������`�����^�R��]X/�Mi6r�6�8��ؙZ2�s�69�vl20��:���UԲ��l�j��[�-t.g���c}�]�-b�7ޞ���n�W^�UID�Y��p4�⋳q��H�x��;�~���O��c�?���
*&���B�H�
/Q`