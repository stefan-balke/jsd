BZh91AY&SY��0 �_�Py����������P�[h$kAA$��M=SSޓQ��zz�5=M= ����Pi�FIP 2  2  �H�h  h      �&M4�dd�т0�F� H� L���T�Й���mF@�����"`�	( 
�A���[�|�Z��4��5�?���]�@�ƅ8��GS)� ��
[f�����_��w��{������+LC��|�ӻ)��	c�3�ۙ
��O7Yݤ��ϕ�m����f��Q�/4�ybH�61\I�&�g>�-.�I$�~7҉�`T�^��i����p�K�Cv�ִ��3&���Xu�s�����(���P�c��u����a�C'RC��F��ʠ�����d��C�'+��i�#����2T�DS�BB��vp_yh��1sU"u�'�d�*�(4��d=����"r�:"Aʄ$9J=*	�`EQ�Atj���[$\*)"��:��9�g&i�k��e�*� p_ �.,�3e�D5�E��𹧓\n��Mh�ֶr�
���j/j�˸�5���m��%��d���4�B�ؑˑ�R�$�k���5��MI�H��I	CI��kj��EEʃ)d��K c@�J��II���뺽e��>���	����{�=�����a�<>(?W��0G:�8|�T1�('����]LI\�O9���0曪' %�%��*�����6�G��rB���82�c�a�yE�L�,��p\`)_�3gITؐ��h��Q&s08.�+!2��{}L��΁*����N��-Ǜq�sPod"(y1��PL��`j���r��"��*��g����χ���_�I@�	ƅ[��_@��f��iq���(K��W�M'��i
�E�%[	�t_|ۂ+��q��d2+��V7E��V���x�H1��.-~x�fHT֢Ҁp��0�m���?1lY� F�	ΐ�:N�&S�����16����&��h�泛Ȑ�`@9h�D�*����Du�B�M��-bT��J
M��J&�������mܐ�������2Fs��N��dUhp�q����S@o+�:�Bā,�bh�Ñ�␬��厃�\1kyP� ��s@�u$@2a��REG��-9�R�8q�1V\\i��X�BjN�<%L$2f�# �j&�(v/��Au��g�Hv�r*�?H���I��8��e��c���Y�so���b��8�Z�{���o4,2.��ܑN$ �u 