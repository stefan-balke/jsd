BZh91AY&SY>�~� �߀Px���������P��@	T�D�ɦF@ � �   9�14L�2da0M4����%2MSOU6�m&A���`�9�14L�2da0M4����$HM54��4��d�4�馧�Ę��!! ,���~����U������Ĝ7�H�hW�M�IȈ@Z /}]Gm|��4��I�����$G����x^�dR���Nʒ�u���sx�v���o$���y�9��#�Z��q"f�f���Ǔ�h(at� �.g�g�=��P�|��`7�/�����RT%�1*{��f�PE�H�΋�Z���#T�sL�ĩ[U��v��0(����&��l�nn��\V�%b�8��#�4b�^�L	�C�U�<|���Į��;xj/%ȵQ5��$!!	]$�P"3kd�|�vb3|Ɯ�ASۑˑ��`!~��T�% �S
J��\ش�C�>b&X^FZ�! ����FTP%�+��� �H��b� \�@�vm�����D$Tm������`E��s�v�K��D�EC�)gچ�-�<8Q�r^=w�	�#�^�/O��~A܋��Ba���F�v
a��H�}1>���]��м����Fl��PL�`h�d���g"
���A�S�$�J���T*l:��vj��P�N��(Z��I��&a�)V=��(p3Ǥ�����4���e9t}#�X=��E�jb��.����3�0h9�醁5�$�GOM}�v�ɑ�P�IMi�;�̢���i3�3�Z>E�X�QƂ�Vƈ�^|a��k�ɵ�LHٸ���Ӽ�b�c�l4�bb#pP`dL54NfaXnz�(ȘG6jH&@�Y�DA�/*�P���7.%h\Q�pz�$D���w�܄�Ю�=�3Y�ց"���D���qA _��%��WJ,�"�h4&W��9�Ą>�+��:;� �2��j���/�.�_��Xm:�g�(�=nH������͚n�U�V�݁��i'P����T�I�MKPb58�--}Ă�u��PEg s#>e.֑���5�ZLY�i#I�@���:��h�E���7��><�6�F�K]�33a	F������"�(HX�[�