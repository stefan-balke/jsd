BZh91AY&SYfR�� �_�Px����������P��@,�ڍ 	IM�4Ƨ�� 3P�4�F40`��`ѐ��&��DA4�=MS�ڍ��  a40`��`ѐ��&��E4�ɦ���)����@��i�<���O|B B* \������,Х��K_�m��D���\e�CGkP���+����3�8A����9q�h[e��#�{�U����$�8�RF�>��\}�����a�β
��R��E��hw�m)V��e��0Z��s"�n TZ���~�k��[4��->́Ƕ�сn���2���U
6���Tӈe֪`�F�-mʦ�i�Fmc��̊h�RE�&*�Լ�i���S
���i�Q},���sf�F�إ-,�s��{^^�<C�{���Q�t&�**>��P���7��m����|<r-�8��X�ބ�(T�6��q�i���彊��"�n�" �H�d�Cb
e$��k>+�m\ה�C~t�,����.��v��G��M�
��#--�n߂���>_d%P�vc�C�FZ�琠��<m��^i�@{
n`LC�,�P[�h�A�����0�����%�l�_1��Iy��׵�1f���*3`m_UiLd��B����<�;N��)K-���N�۳PuY��1=���PԚ�i('X�g�)�fk��8ϰ��Xg��qL��@L�aD�y:4H��uA���c<T���l!u�����N�,ɒ2���j	U��S�pX���[G�yK��Y0�H%�y�U)OV�hүbF�nA��v���S������Ձa�	��'3����į&�H	ة�����ACiH�`&��q҅KD4@{
$Jl`�7j��	厴��� ���ua�y������������XЙWA���!�{G@1�9�7 �)�u+J�'Q`s����C�8p*rDW���Pf[w�$�\��\��MC��H(]nD�r2��jH3,+"�
��UH�`�<u��=x�M��&Akb��b��j�H��A�o���3UWg�31$�`��]y궯�]��BA�KG�