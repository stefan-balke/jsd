BZh91AY&SY�	�p k_�Py����������P~;g�ΠQր	E2L�������#@ 4��Jh@��h4��d�    	L�(�        i��ɂ0�#M1L� $H�d�L MM�5=MS�h 6�z��ć�@�@�@����g�B
�)&�4$����ہyM$��,�GkRrQ	�JAs��t���ϏE���>��<V�^�-�Q#���X�Y�ȵ[i0�%7�}�h�%�M�?0��3�3�X��<Vۉ�M�:̻
�Z�aY��δ<γHBwf�SHC�dsa� W#�5_����#��eրi��=hq��Q�Ձ�㏛9B�#�IV�Aܤ-��Z73`�f*�vg2���� xK��4Lp�Ƥb5�m��[Ve�%4Z����J������EI�!�f��4hk��0Ľ�����L�r �_*�hW1iD���V�D�v���&&���a��i��,k�tcB���*��/S��ۼn8�$!,�I@�3b�u�*H��r�!U�H���*��hM�Q�]�%m&�Z��j�50�6�& �E��2�� ��ll� Hl�a/�������iü`��0������a�iH�wG	'Թx1xRZ3Z�0L�|�I��<\8E�*��TèMž���[���7��6�+��?���jW����v/��P'�`5AF DT����)��Z-SM��5�*3���|,�4C4�ugs ����I<(�r]LS21rw��A�����|�5A2�mM-�%�`��JK�x���C����uw�P!�8ġ�HX+�?0��A��b�(
�w�w�Lg��hnjf�E"H�dt�W��� �DkD!͍����iHN�M�P)6�ph$�rr�&U�� �:���ֹ�kC2�HZ6 ;�'8��r��@����Eraq��B��� � ���$(1Vꂑ������BХ��XĩE:��*Œ�<�1]��r :Mɠ)8�B TCMr���;D�	a����@�\V�u�Hj+�z��bB��h�a���,�<UŎ��d�ɺ���FӢn�2C����RE�`,v��5���U�V��z�h7䙐��jN��
 *e��!��C �5�[����_bAk]M�Xa"UA��4x)v4��KI��A���4�"ƹ��a2h��kn�f�6��UKZ�ٚ�P��_�����"�(HX� 