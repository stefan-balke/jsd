BZh91AY&SY]��#  ߀Px���������P�q�w �rwj4�Rh)�=C@�OPz���h)�i�*~��      S$ԛL���A�
C  2�`LM&L�LM2100IS	��� ji?T��Aa��M�$��$�$dBB���ګ��{��%Ԇ!)z��~���=��xE�2�D���v��Go^�U��|�ݬ��-�܇�p»҉��P�ch�f��J�!N�Fr�Z)B��Tډ��٧!v��(�f����m�4�&�r��^c�$�U�6Y�z��u�Mc 3ۻI3Dk'+?rjy�\Fnl��p~��BJ�j�m/Z&�������m>
(Z��$Z.�f�n��,\�F�Y�N�B�1�Aa�fM����VΑ��V�T�B�j�i�aMz%6�eR#%>Kf2�+),���C�.!إtφw��<�l�Z�Ќ���6�,�M�.9�Ҭb��d��j�f��1d�R���*�4�p�84	6s���寭Z�cPZrEAl��fQG�\B�m����"�0���>"��6x��N!	K}$�P"c8�'wpyf#��,��U�H���+Q�1"n3%E!
8sbd$J)i�!��&.�*j �L���l���r��ẚԑJU!�R�b�z���|3G�1� pyL��?{Lu�s�Jګ�=��X�S�	h	)�4�rB��Ew'¨�X�/��o=?�֤����Zu��ȟY����=_��m��ϐ�>%B~��c���^���O4����8�{g�|��	�SN�'����9���|uS����)�s�щR)jrd}]�8��+���z.��8�]%�f8�[\aRgr��%�6�Z�H�Hk^IR�M���&��#�n�	��as<a���=K(B³�0*��R�1#�X@<m���><e	��y�^;�>9�Ϲ���"�@� �*�rJ�di��`G�5���c�X�����,[|��7+�<��׶*:g
�d�V��x�B���ү�Tr���88�t�(q`�D��a�����Ł�k�� ���[:��|�X�J�L�ܦJ�3e����H��-bۻ��ˬJ�(O���|�!����c��}\凛�gob�0�8<p�I֨�����拢W�p�Ey�(���	�Č=�fƏ��<ە=2UJ�)�޺�&Uh���&��j�N]��L��5�:Z�v�fb^�m�e	�m�S��o7*Z��ri��sM#���\%�p�����>���RTO�g���l��E�9ͬ���gv�?wRo��i�|��`܆@�0ѹ����ܑN$gm�