BZh91AY&SY�� T_�Px���������P~��d"�:Q�A��D�SFOQ6��z��0A� �& �ЀR�SF����  �  �&�4ш�z� 4�� �=M4�sbh0�2d��`�i���!�H��F�e=e5OS�2z)�=L�F� z�Hi$B��@�@�?/�r6��,Z���XI��8~pm�ـ%�hUeX@�;ڔ���@j~�:aյ�;s��8��4_M2��w�`�9u��m�P�~�����!�?v���..�qg6��,\�
xWZ��]�m:q+[�F/�F'{�b@�����������IP����O)7��>僌I�}��or��fd-��K���TUKfڊk2�~�5|.�	�L��4�+a����X��:�,��h�A^Y�t3��)N)D`�QZH�Hl�̶(�ۭd�t��e���)k�kH\4�0a�m]ب��i�g���|�SA�-�]J�i�k7��61�-��CIB���8�-|$r�I;NJ%J$�����@1�i�61�X�)��b�X�c���e�1 ��  :l�n2Ck�I)�T2�t3�,�' *�>3����
��k�֔<��?X�sB(�<�����3�{�-$���d���k^��I%���zu�p���-�1/�!и�~Wt
a��ف��=�nf��1줺u"�-b^%�m��:,�l}+��
��o(]��[�OmVY[isc-idvb\U�72B\�ƍQ&P[���С���2׊�9Y�֤83��Ľj�@�	�:�
����h>�[��#Al&'�x���J�1.2�%�I؎]vx�p&FV!���O�-��L��4k�l�
����⸄M�
@P(`O'�bdZ���f��0���A/gxe����e@�o/*K1X06����B�n�NSh�	j�@�=�PbX��bBB0=�VH�dvo�0Dh�y�I� #�km��4=Z!=��%�q	��T�<�b=v��Ӂ̸$���#ՠ��Y�	��v�I$�X��2�u�p�&�����eNәh\/ai�eB�m9 g���8D��*_�hZ3[c��t�7^�P��K�]�5�@�ḽ^�W��Y���Y �F��RZ��%
����Y�4�<�Ζ�H�}d�Y�L��S)�Y`Ip����Sk�pV[��f#A�`е^w�O�]��B@^�/�