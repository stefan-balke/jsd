BZh91AY&SY�J`6 z_�Px���������P~�@�hh���Q��442 �  �4`�1 �&	�!��L����j�4��=OS�j �M2 �m h9�#� �&���0F&(S& 	����6���C  yOI�.$�=��SI�
���9F��A��CIX���{�ۂ��IhhY�M&���f@������u�������|+A��S(��'�p߾ai�hӦ6��Y`F�},����r�����Pe�C���H�'ytu��U$�qu�h�w{�IU��R,�����V�x����. �Lz�{8��F���y���Z�2��J��tQh�*|K$X�܈0��"�y2�i�XbC
C�dbDav��f�/R�&ê������b�ϵZ�#-��^��b�#&KlG�5��L����nn�-G}v�F6�QЫ)�5��2��QnU��(�G/�˴Ͷ;l�(��c�4b��������t��lc|���C@B.���ZK�9P�玉R�2\mbF�H�	�e��B���A�i�.�(da���k��b0M�h��+�E��a�>��am���@�����J	j�^��B�	=�`ax]�)��H��l��彽��Хċ�9�U|�سB	��!�>��˫������A �o��vqH;��\r�`y-��Nu�2ͩ/[�D��1f��0�����9H�c#9ˇ��d!�g��|�
�3��XΜ�ō@��"dw��LL6�nL�Q��F�As�2^,��%�F�
��{`!��3�0�;��=�5b�*B�L�i���<qL4CA��7Q;��Z6$Ȑ4؆�JhZ_v�dְ�H������ڃ/A]�|@޴�2�]!p�*R��5��*��-[ =��9�u�a�ai�1���%�$��R3� ܳJ0ĒIru�Ab��$$#A��a�2��"#F�`A,�f"���=9��p7
@2��zO���ix�>ϙ�D��5�Op�<">��4&Oy��@>`/�x1�?`����z�V�8�@�T���w g.�$�D�Hp�j�C��f�|�
�E.KEy�dK	P$��[��c�Bs*�A�a�2�*D,�`u��&���ŤH�_��^ji1���k@,4+J �@ײ��י�N����h4Fe8����)�JS�