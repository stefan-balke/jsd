BZh91AY&SYz}�v �߀Px����������`��s �4� !(�S�m53J�44�   ��%4�@� �   �0L@0	�h�h`ba�����d���    �0L@0	�h�h`b`�"#&�LI�a4h�6��OI�5�V0J���R�"Y
��5]�'�heQ.T)z���U�G��J�fS:,����֩#;X�^]��y/G���-�7�����x�1�331�0��d�S���/��qhĈTWI$@M-��+��T��&�TF�I��#��D���ݒ�B	7�tYM#"ȋdI�*�	.4
�ũp9Fz�h�"fhG�N>j\��eUU2�y��6]��g<I(�i��W��Q�W�lg�mI��ExO:�%���@��AA����xw�`�
O�����k��U�������[l͌�CzJ��T�� ���DMY�&@� �c��ő�vP��΢Q�!QQT�4찯=em,6]�p#  ��5�
l����9Y��}L	R�D6E,)Y.���1��T���gC�˧h�l�Ch��Zb��iȫV�4�ɘq��i�E6��M!y�f��!b�Zj��D�)�e�KSVBM
�;@`E�2�|ux�N���Ң,l��v�K�T���K[L�"�`b�j%���O�@�At D(��Xh��%�*80&9jT"��S�)�E�UZs)�4L�
)���� �.��A-V�S,P:��D�2�(���\R�������gu˔Z�k]o�R�UF��[]�y��e!��{#K��@w��zW�|eÆ���ϮA�r�\^>/W8�l
�#۹䅂�[w.A�AX�7
��G��K�=T��{n���bG�;��^�������#Gr��,n86=���N<�)��KB��}u��S�\�ژ��H틮m��灔��C|�g%�7��g�]��V�K喍;��JV�GCǣZ���}-�ߪ��b�c$r�r�	K�����Un&���~�p���W"��  ��nb��fe�S������ojtLR�K�������a�,Q#��S	�/'�8����8v.0�芉K\�Z��z\&A��<�)����=����M;'
�b�W�m}:M��Ye���RsM��tu>�h��1�W�^��M/I��n���3eH��+Ua�
ؼ�5,,]ۺYLV9૭e�G�[�e##Q�t�h��	��&)z��٤�aK,[[���q�[��$x9&�͒K*G����ys8M�a��Y����I���b��z�qY���;Ďըs��YE�.$�s`�s�,����47�i�d���)˒�R�������b����c%8�vnL�&Z��I�����da/Zuv�$d�u�Z�u66�,�����ɣNk��xUc}ͳnp���Lz�F�untԔO�g.N����f�R7^,�����]T�uLs�G��:��EDհ����)����