BZh91AY&SYs� �߀Px���������P�{����F�j�j4�1=&�L�#F i�h� $�'�1'�M4d�4a��!!
#&�1���&�� 240&&�	�&L�&	����LL��
���S�S��6��hh4�G��Y! �,�@��=㣨���
�"�e5>��q��#A�d3&���PH�2�4|;�����v�����vi�O����T���tV��P�k���lt7أ��ۑQ�6h01�/ �9�d�JMgyLg�#J�h3� D�!#ޒDA�f���>�/��&�1��9���#E������:��eR��QN2�����՚�Y��mf.X+��h�0f,q>�Eɠ�`L��w3,�����j��p�YX�Gb#24��*_�X^C��٨��8�lczm���!��5x�Irpʅ'y�T�K�a�mI�v���WXw�-wZ���T-�PP0�p�}�1��k�����9sː��Ĩ�@㯗S/ �"EVhր�u�G��y����׶��Q�ww�VG�3LvL���ۿ_q�'��a�-�b�@b����~�L<A��%��q��V�I:S\��etS"�ύ�f,��b	��l(��A���I�J��ܪZՆgm�C��5�B]����N,ژ9�5tR��X�g]oC��E����48ȧa`W��`bv�a�Zd�(
�:��L�L�H3$��#�G_]z��9�%��4VSB��5�(��*g���w���XA�ķ_V�`��f���0�yV��ݱ-- �]��x 4r+�>m�t����[�F$�K	��
�s�uRq�D#G-J��|K�1!t�\5�a��*9̩4CEB�D��߷/V�'��u��@C���#�q`}ZM� t��H�n=[VE�hj+��Na$�1M���LTA���T�Gad�:��� x̙�À�e"C��������o�U�V��v�}�,'P���w��t� �5,��[J���A �������H�P@d�*si�=��MI_a�h`kR,5͗��7o����ک�6��?k22!c�v��E?�w$S�	1Q�