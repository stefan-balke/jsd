BZh91AY&SY| �߀Px����������P�v���c\�@(��i2�S��=MH =M@4 �ML�4� �    Jz��)��OP4�@  `�1 �&	�!��L���i3CR=	��?PM4ѐ��jyL	�O0�B($�w�)�����U�Р������  �_C�ud�����`�a	�A(L��l`J�8�n�&�7=��5�'`��Fɦ���pd�j�'���p<P����E]��S�;�1�;�d�ǻ�Z�eFXP�s�^A�s5KX8' e����A�b�z�%a���U��v1��v�&X?Z���}W,�t[��y4��m|���*((�ϙ�Az�
�#�MH�}Ü��J�@��ɡ��:��С�7 �t�j�KOe䖋$TcX��J��\Q������&3i�X���
��\��M�R�IX����/�C��MV.ld��\�
b�SCu#��t�*V�S7��!C4c�����EI�X�yvqAr vp�%$�]���UjIڢ��ES�-s{��a��:b��.ꪰ D�qX���~����I@7�*&����[Р�0~*�E3$X���j�/ �,H��˕�p��/RPIl�((b�$�h�TH|�����d}��6�w(h0=�����_8ф8��V�!��Y!�$z�
CJ�.I�w<=��b�5F��!�UV;(���6 ��t��{þ=����I����~�ݖ���nB��@>K�P�R���%APS֒;�0dwT+�b�	{	���TD3a�P��d|�x$�,�J���-	���y/��A�!C��f� e�����B5|R��U!�9u[�r>��浢�(�8�(��~�� ��k7-5�
���hz?��릻HH���A��B�E�#��^����mȄh��w��l��$��������uS9����Ε*�|W~��z��<����z�p$6�Ir9��ħh��Ph���4���*D�KA9�°���HH/P�:�PX��,4L��rx��VI�1"�ju()4T=E�M�o�6�}�Omv$�����iB��xzh�����-�<^�2<��5��>��4&W��3	 ��I4pK ����$k	�@�߭^Zv�����]xTm: fy��Ɣ�ÜK�PzRվ3(3n��
������a:�ԝ���I/���@�y�d����~,[���%T$�c�R�i�=ؙ4���H��d���a�`U2C ��<_#���Z]����0hXP��rE8P�|