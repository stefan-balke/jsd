BZh91AY&SYկ�	 �_�Px���������P�wv�q8�h$p�4���Hڦ��   �@4	�*j �  @  $$MS�S����j�?T  ���b�LFCC �#I D�!�=21=DzG��44�&��Eo���0�eY
��~��Ƈ��Ƣ](/B�T��������gTL&a�G�T�1,�4}���w��??|���3�I�����_;��tٙA�&çSl/#�G�fg0�TJ\t� ��nSv�7&Ν���^��ܽuߥ��S��`$͖e��LL���0ϒ֯�c��_���1�]_Wxs��ݠ�딥�K:"�v��j^�:'J��^�����b�t�6z�����jbXtÛPn��5v�1FL�=��W֕�\�ɕXfl,��1�Fۆ�����&X�֊����$�N��J�T���Q�&ּ�/83S��7R�I�
�$��	(KJ���,!-�
s[���҈ӿC49�61��m���B^���>K���T)��Q*Q%�]�fz�j��҅�M�,P�6�#rF�Q0�I�.2�J-�#]�_f	���ů��M��<�\��w�Qcw�=>^���X0��8�m%��C���L�xN!�S5��+=ҭ�b`zb؃sL�Za��e���>�����8~'�oY�F~E!���f�mw6�ڗ��-7�|�CoL�)��'˂|�R�I;дk�+぀�=Y籠&Fz����d!�1�{\+,���ɶ�lu�9ZY���x������S�T��DX�/�b��jW6y���w������V��Ѵ��ʯH�W>~S���^�0]�����z����y�_;GFQ�V>�6�����G2Z2�����Ʉ�5K�7AH�Wv�K1`_����2UP�X.F?h�,��<T�f��M��C���L{�6�q<��L�o�j^hi�0����uV��̲ � (��PE�;�,HHFG�r�218�2���C,�.���ȋ_KX�\zӯtJ��c��B`)�ݩ%�#�w~G�����Xt�,�o�Rjp�]��D�N��d�B�CL*:�Q�Ýe���3�u�[�Ρ�ɑ��U*�S.(c.�(|��Gd�`g��(�������̾ʞ�x�dkC!��oZ�5KC{�~,ˌ�T;x��c
9+�_��u�SeIR=K4���,6��f١�5�o�7o�῎�{��g�)��hs(28�r)�.�p�!�_^