BZh91AY&SY>�5? q߀Px���������`?z��18�@J���4�z�4  �   ��)`	�   4ØA�ɓ&F�L�LBF�5I��i�i�����~�� �jz�9�14L�2da0M4����$A &�$2)�dmM �F4'���HWY�c	3�B�/��U�	/� ��CH0 Mw��6໰ �*&jgE�Q�R�Z��&v����<:���QN��Gr�gR��5J���P^�V0*�3�����k�TT�������dK�:�LH�?�g��zӞ��d�m
�m��Y�V���i�k��n��捳�k��$!���1�I�����4B��N�c����1��:ϼ��X�i������Q˜�^:���K&r���UɤWwNJwF�١��0����u�F�kF���lc�cɉ[�̍%��;X�.)��v���أ)��F�]�,l��sB�v��̐�k�8�&L��m��#�E�a*�f�)�i��,�jj�F��͎&n[�J�����9�^�^[���8%��G*R��L^Z�0!P�*+%,��J]�@A��0��\M���%�n��HPP-���Hr!�^�JL�`Z�	Tz��<cc���CHC��:�礹|r�P'��T�U�f�	�Bc0S�����e橍�27݂Њ11�64�1�u��FdD1�#^Sw��I�wM��잝o�5ӏ7��46?x槡"،��'*X{���� �������k�u�%t��,.�M)��
BU&|.0ZA����^s����i֤�hX�k{k�wk�L������=d�꟢�CGY'��Fi'փ�)��bb��C���ؙ�2�;!�Nē��Uޚ�.�h�w=���YƖ�W��n�1%1�ڠu&����5�f�'k<����49֟5����Q%[{�3/r����z{���)s%��Y���w�RE�+�b��(��e���,�Tc|"q�lg#l��/��{�9�V����H4��ŋkqW�ƥo�,��9�Fɶ��ݗDs�*=,����q5<L��40�L�706�L0p2�V:1S��܀@�����y��BB4/��H�ll����"4Xz[
Q\��ˤJ�ù��
m~ݰ]H����mrl,=M��oz9ϧz��D�^�����
��Q�)F�o$�	��if�{Jx�l0UJ�
v�ԤƭV�k�����)��=���-g]H��ٰ��^����MWYe��l�j��6'\Z4�\�5ō���vP����/��u�s�II>=^.&��7|��&�ŝ:�s��]T�]&:3���P⢢i�[e���H�
ۆ��