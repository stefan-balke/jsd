BZh91AY&SY�ܥ; �_�Px���������`�z�g A� 4��!O'�<������� �S���4�     9�14L�2da0M4����%=$D�4 �     ���a2dɑ��4�# C � A1&M4)����4 ���1&!x�$��$� �@����r5�AF��T��-��_\+�*�^4+�@��Ԝ�Bh���tpϥ=�2�=E�Z���2��K~S�m��!�p2wR'�w�@��*�y�
|Z�RCnf�]9�9�q*R/�J��0���K���<� ?Ojb	8��m�	�#6fj���$��ʄ�����t���e}(V�3A� �J �Sxg)K��mΣ��1 �������AnvBd��<J����y��sH�9�X����*J^�O�N�I�P� �K���B�̹<Bt �U�񑀈�"u62�D3�
ȗ��D���9��ɰ�&�ki�cF9�̒��ժL���:���uix��f�A̡!�*���=V��L�Q��"�r���W&h���r����m���V�
(M��_loT���ڊ�(:!ښ�$`+pQHl�yyk4�H %��+&uO�@`E*l�$�j�
F-�����q��w�s��w�o:0i��ie�1͊�����7�D^"��%PB������xzde��ݒ�cP�+�ۋ`���_�A��dj�ݬ�Q!������Et�\	���]1��F��ɾ�KJU[�w�����<[���Os� �t�1�Cs16h_ٞ�[�I)�W��䂏�����4�I)~\|CBU(�����G�!i%mrK�"�������]�x���.b�����@�v?f���x�!r�1�������j
�by�Fm>t*&�U706����Hd3a@��E�RO:�[]�K�.#�c�Pld"�����P(�o`s&��"`�΃�Хb=��]Hp3�yc%z$�i!ƅm�`�p��fu��CYx� �.����Mz����ĉ��h�:�W����$z�;��i���n�pf�bL�a�?j��l�S#jsa��Р "��hb=u�{�7!�%�-��Bwq����X����Q�q=�V&4)̃XVM�I�3&X����E�9�`����&j���z'0e�9�*4CDʇ�	 �� "�;�A�xoB{k�<��(4>�=d���ං��a�b��2����A�p�0�	�Ѕ�GH@Çh:�E�q�v��]�T0
�49yI@�4�8D��:�yQ�8��a�7�b�3}�.'`���R�AS��d�F�⁾���H-a��),�Q@h�K�K��g��374��a�`^��
E���ZI~����e�T�+L$��Ҥ@�PT݂M��.�p�!��Jv