BZh91AY&SY�W�E �߀Px����������`	��h  �ϽWT�:��ҙL�Q��O��CLe@�  ��h	")�B2h�b0��4ɀh	�2d�b`ɂd ф``iH���i�@d�   � �R��<�&�mF@@ d �M �"L(�'�d 542  %�$IcE	�T2�V�Q�B1q��� �a��`C ����%hqd@�P�iD,�0�f1Yl�;��ѷ�'X���).-�Xx��C�<D]�
���ԣҏEB�Hx��!�DA
"�!�R���r.�?�ہp-Ej��$��;�`��8��*�1e*Ҏ��pv&f������h#��O�/�������,)Y��sK&��ܒa�Ț���i�!Kr3b�dQ	�^RU	�C�31 �5�G^wo������ڪ[��w�<�|�q�潷&@�M���9PwU�m�Y[P���#o-5�8.$��!B����p$C���I҇wPA(�N�7��>,gq��O�?�"�>�שn�  �< ^!�q-qʙ��I@����	�c+�E�Jb�r,�Q7�T���C:��l> W܉����q��C1,;d�d� ��°����㩉�"]�$ �����M?~���@=>m^ˇvQ��C�jp�x  �9�9��C�;-��xY,0I]�yp`�{�8��\8��v��gzB��GT�f���@�l�(�@9R��l+k�D�s&$EZ��� ��$p�9CD�j�T�q�KY`$'ꝥ�!���n��`];Nڜ7�N�ڨ8P�Grn�\��^H|�r���$��uG43-gb��\�!wf_��6���pM�kw/�]i�Y�G5P�Z^,%&�\T�ڪC#h���L㢋f@�0AO�w���/.�W�Pa8P��b��M�y�TT]�Ff�xL4٘���vB����DT�u�u̮�=����	<\6J���D���̸Jrm���{+*/P���}��K���S�d8r�Gg�:�����)9�t�HA�y���Ӻ�x����&dq`O9��p?��N5#!
�Bx�W9f-G��!DQ���@��s#��<��+qL;��qp[�Y�,��VQ�9ұb�S��(��,�X�b�A�E�,��\bR�8�
(�2�DH�#1J5��X�u�1�Y�%2Չ��!Y�zn���I�����/������a~1��q��#���cl����(��z2��t��0?XT1��|��M��;������$���%�V}I$�Q��)�� ��K>�d�n�l>�2X�t<�wk��zdt��,=��;d^WqVH��9��X4 ���UE-M�~G��K,�4zd���e�V��d���H��׸:2��as85���)��T��K/�E5[�/����olr �8��jj�	(�UTd nٜ��32�+�6�ӧ��hn��+�����݆�b�N��\)L'�x��<>�gK�1pɄ�e6%ǖd�0��nbF�":�d�/�k�l!4tN�H,U��\��5+v9e����6ch$�q!>_3�*:�����߉��lf�z*k���Z��V��$�,,]պY;X���b��e�A����##��t�&����a��I���BZ�vڮ��b��@��i���%������h>}Ι�,;9���=&�Wn
��D�^k�f�BYn��F��v=HM�� ��t��hx�V��1�Ѭ�U+T)Ϛ�R����-*lA��nlT���beh�I�j�M�yݛ	���i��ĄɎ�Yk8���
�K����ѫ5��P�nJwWU�� �34�V�3�&b�K;M(��g/����ٸ�L�or�0`�b!�]e<�x�I\ !�J?�ܑN$3��Q@