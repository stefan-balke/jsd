BZh91AY&SYA+�J �߀Px����������P�	��g�YFE�BEdѣ)�Fehhhz@�4��d��  h      ��T�*z�j?"1F��?SP�h�Ph8ɓ&# &L �# C T��	��D�O�4򆁠@46�ad�����2/{HT ��t�r��$�$25���F����A�dF���6�T�ID3>=�k���Ѻz��]s�ɕw/�1�yq�"C�/���m���ZDyS��v�9a=#�4�m��'�ʊ�"��l-��jw�ci�J��dGF�T���BJ��-`�_����\�8��㻼�adHi�s~=a��#E��E޵p��1���T����T�x�:3;�٦(Z�>�z�P��<ߦ|^���
a��!�ҙi�������֝�	I�`4����-[Q�%P5*�@Ut*�ܦX� e��-���D�4^��e(0�$�\�� Q��X�y�!y�nU����d�h�4U]�7��2Rȩa�`ƛs�M4fy�x֦��u�9��61�V�m���C��G�:�\:H�B��e�Z�&5
 څ�0C����ԍ��w�L԰�G\j���"��V�nbЛ��6��}|���E��G�xg�:=}?{M>#I��t��f���Qq���v<xO��J��9���A�����g�h�RG�u{۹�~��o1̙��"����1�ݙ���nӹ/<
Z\?���#d�T˔���OJEF�o���
��(�ũ����dE;�'udªR���WD�G�����V����q.t�� �t`ֲ��3og�C��ۊ,�aA���4�ޱ͘˚�a��9���f�zX��/�=OI���n�t�I_^�º;2���~S7��1�)A�HY?	,��K���ge�X�~��w�`��>���bŴ��m�{����S]��M�rH��<Gc:���7�hh6jf]�LT5�5Q/����W�B��0�i, Q��Ab��$$#���\5
,����b���(>� )fH&����%o��rGs�0��.R=�u�Fc����Xy��%�G�7+�ڨ���]fK���UR�vs�H�_"�^�����:��p�N��p��c�a�U��D�j�,�;+q�"P�aR��f�B�Y��4�-��3.2�R6��� 䁆�Υ��.�|��	�������2n��ؓe�hp�c�㚪{&W�̋� �`ЬW���rE8P�A+�J