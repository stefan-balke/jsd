BZh91AY&SYn+�� �߀Px����������`Q���w��� xJ$ʞ��hSy"i� 4@�=4�H�4m@ �F@  ���#@�����@  %=$��@  h4    8ɓ&# &L �# C � BM115M�a4OCS@��L��H{�	@��$����G#8��hR4��_��n�4 ��Y�h�jR!�	
�{��ݾ�w�ߖ�<���=_Z{֓�KT���)�Z�+JT$�T�̜��ʍA)I(@�L�<�ţ����8>W<����JCn#C)ɖ4�yg9oyDQ"��A��.�a� L<c�0��:�]g�np|��������Q�/9<�>b��e)FD�.P3b%�Js�A����V�)D��S�bL��g��(���o�/ë���0�
�
-0�\!ȡ��=,�v�#=��9Z)�73]��laˎQ-���fV��OQK����`c���X�H�Q��C���w"�*�Ź���e�4���S
���V�&��h����U˖�C6��sts�^ɢ�֬��5H�k]��S�EƧ�.W�wV"[+l��f����8@W�g�9�EL*���#�^3+�ҍ��MV��2�k�M����(��l�ȭ�n`4H6ɰ��,7. J����T 
�)D��vkV�6�޸��E�(?!�S,]�<hG��5�Ye���:�B��c��ǘ,��D7Q�f�?N��tU�kѷv��Y�x�XMÂa�ڨ���%�6KM�9�F�RCN�Z��V���(l�;1���v�in��cy,de�gS^�q��ǚ!�2r�i�9�7;�7�M-���i�v�緽K�.��x�ɩn�r���b"�1�s$����e�01-Yx���^F��@2b��-�[�<6�C,��î�W���Ex��ЅB�9[�ϲ�7�˅�NS~�r��Y�@Z��F1j1#K�p���%�.Q��@S	y�������iZU���R4D$ H]�W],j!�AP�vXX!�nM-$��!����M���u��[<�N��hyu<��U��/s�</Yp3w�P}Q ���j�VTBN�m�Ȧ�JDCBR"gHU�4 M.���Gxn9�t��p}#�i+��H���A�g\���@`S="#e�|�z��]��!w$�#&l>T
$ͬK��i�d3P��k ����$�J�����s�}�LŚ�������[ڠ�( ��[���)XR�y/k>�Mtt4+��@�bCchClb����`�H��be��������%�w��L���i8p�����F�#����״��!����Ew�trZF��X~z��'�d�]�r���|Q��`<��-ly�!�BƐ -<�=�'X
y��r��@���m���L3���d������ $s�D�d���D�_�H�^&��Z�5:��*��B"l`�d��'�ɥ GA��f�:AH�����K: ��j6A�X�{(>!�4&[��o!󁐓F �Νi2	�L��^X�yK��������7n!��D"c���%���Xf�kha�7`1��,N�5'~�$���A�g3�a���P7T��Xb\[��V3,���de�R󴌾�fF�� ��m�j�bR,kXIb��6� ���mxʗ]w�̆��`Зcg�.�p� �W�