BZh91AY&SYK0' �߀Px���������P�צ!�;��v$a(��M������ 0# h�SI�$��4����    HIj��=FOA@�=@ 5 ���&L�20�&�db``
�@��4�BmQ��Q�=L��#&�C)���@���K��Ǽu�A��/hT4� �k�E�{�$gJ��Sm|���j95�ǯO���`��L�t�r�o[�[8����)�*Y�߹���G�?[���`39�v�c��)�yp&UUM��yNq0�gL�"�������=�J���X�V(0cͧ��vDg��M��YI���@��Y۠T�{h9�6�2���ڱ䰯��R&��AQґ�HMf�|A�:�e���~j4͂�����b�+R��E
	���	�R��_gsw�!��T%P�u��j���m��C��k���G*�ߢT�K��q|�7W��)�6�#rF�I�A��{�z((F��g�l43tƛ��&���3a���\���v��Tll�<`DRc��������!J �Nc��r�I?�୍U�ҧ���6� i
�$ꎯ��S�:���H(b^�ާkf����%H�Dc`�ǖ�ޘ�%w4Dx޶#�x��n|�-D�H�+LBb��a��>��s$)Z��WA�8s��9�C�%8��M\�]��M
�XХ��W�k8��D�>��#?YD$�kX�ȸ��>��������b�P�Wc����c�I#��j���T&j֛�!uq���AP����[���%+�D�=+��՟q��f�F}1�
_9��m�ߺ1��-�=]��L<�|��2���^ש�\p.H�Y�ºؖ�f�u�ȲHĀ@�^�PX���bBB4zǡ,Ć!�ARt�P�x���[��"r�`��V%���
��Cʿ�ߜ��pj(8�Q����N��%����\�	�	�\�={�%en�cB�'��27ZC`�$�,隡�@��!��F6t�R�87k��v+��&�[P�j,g�`�����cIzb�pXsػ>eE�$䲬(�	5O|W�byN��"Qޣ�[�dh�����/[j�9����ǃ�Yvot�6����h��.�p� �`N