BZh91AY&SY�tVx )_�Py���������P�+����T	M	�MOM&��F�SOS��fQ�4�4��i���&�5OH2�F�  hhMDDH  �    ��2b10d�2 h�00	14�L�OS4H�(@� z�d��P �
�P4���������P4a,B��E���&ih��6�&�j�P�*�j�����wr�螢r�o�8���}��љ�S ���$G�ʋ�l�̰ӳk�.l$�Sh��
"*"�+B���_�-���ŊE���:d��-G[M�yL�j�������_�ǋ�Ā��H�:�`��c�}���X=�ܒԩ���f	����c���bUbh�E[!0�2Z���΍EY�3ZP�V�4���ZgS���<,�"i�lټ�PH:����B�J�D\&-���)�V*�k"�����Z�R�s�|B[E��TA0V��d�{�Yi�v���킷v��A �5ݞ`�9%V��Z��Ic6�\��V��Q����:D��ɲ(�T��Q��`�Y�_[�D�T�wSf�|��sED^��BJ(��3�������.�n��d��Ҳ,q!Eh)KTS���1��Ⲷ^�٣�Q����KA��Q��XX!L�髚C�[[k�`�tÞ���4d�L�Ʈp�:;qn�o�@�"c�K��e}v��i�1�
���쒡�������z�U�R��%4`�.3�.�"��0Œa�]O}KWH���T�!>�`@-
�S��Wp�I`dW��+�+��o�
}�2�[�H�@kH[�s8O	����T�!$�C��j\<�(q����3-�.V��
�CB�xl��5,�P�K�6���,ؗ$�C9��5|R��R=l�\�g�б���Zi4�m �"�-����?X�aA��A�PP%�|��yS^���+�4J�/H�dt��6�&A��h�������I\)���pe[��0c�)��azB«�JW���z�Z��7��������!v��P/9�:���P�i�,K0ULJs1
�s�r�D�# ���Z�	�)���;��o`��Hd$��xE�Ir��D��*��l�����x�B{i�!w�F m;�F"�D5�'(�5�������@���2���0� J�9�G0cz=[���S<�W4�ypz@����A�9�g$�M*X��A���KO�Xf��qa�8�##��X�BjN��HU;�&H� �b�#P�2�C�I_��Q@д�H) ak֦��,���p��K�k"GC`\�څ"��yQ,��8g�p�����-�ɜd �0hW�u�����)�K���