BZh91AY&SYZk�8 �_�Px���������`�k�wt��4B�8Jj�O&$�2 ���Ѡ���M	��H4   h �A�ɓ&F�L�LB!M��<����24h����9�14L�2da0M4����$PF�i�?�S�O��z�Q�����yN�!�"A �����G#��2��)4"�!�׸�-�촐��4�h�ڪQ�Z�6gGY��wt��Qx����.��v�r�l3j��k8��j{)����ud������cm��v�g\���H6�ۑ~�fj��g͘g�%Ha�/!���.06�ܡ,����b�pj{H/Z��4��Xݱ��,R̔<�o�t���Ϛٮu�G�-���$�	ة0�&������>��c/�|P�x:є��׵˛Edlx*��<{s[` "6�G�+V��q��!��1p]��R��I�s<*��Ƥ���
�1:�l��uP(� ˮ�q"��a��K4Xް�"��6Lb�v�r^m�mT���%*5�:�W��T4�dѵ�a9fPAK�Yai+c^��La��Pif4�̭H���b��YUk����jR0�f6�,*�X�
a��mb�$T���p�͜���,�L �\*P.�(�ݷ�3j�d�!���J����0f��z��p���P���7��m�1�:~��z��;/�7���ƅ���Y��Y��;de6H��d�ԦG��Gݖ��L������B8�5TBB)p[�����T�"��
��T�d�� �6���_�/e��8�KggU�Q�FR�ʽ��j�pq3����pTgӞC	�W�z�7�.��D�`x��{sb43�y�s�Y��Pcn���إ�d�Q@����tڻ����J�c@��A���z1$ü/�%�j漃�e�	/N��G�z"�a�ʁ!3�����b��@�3Y@��[ @��r��&1�wŖ6=4.c���oQC�ȉ��|BhL��{A�4��"$dh�`�Rs3D�amȄFy�g(�3��m���L�8���W����ݟQ�-3�*b�xԗi�w�wʘbem3�]��ƨ��Ohfؑ��&D�T4R2B��ͽ֤^��8�3�ݬ4{����ߚՋ�@!������׆�v�z��
�n@�]���'2�[a�a��.(YN�\P-bR��[w�u6,� ��X`��("���:$#�	�Yg@���h�)�A�*��k���/��#Q�܄�Sb]��"h���$�v�GRXn�1:Vw@�X��\��5	��s8H�h	f�&�@�,���F���zVr��2���ZӴ��(��)�P���Z<����A�6���F(H�9�E��X=��.-A�T�7���
�h]D�l�0�(�jx��i����&�� eȖ�����2e�,���|�W6�d�*W�o�cA�����Id����"�(H-5�� 