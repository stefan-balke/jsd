BZh91AY&SY�1 7_�Px���������P8^΢8��:BP���)�4 �i��M@)�&P� �     		�F���hh4 � �A�ɓ&F�L�LE&S�<�����z���Cɨ���yN�a�D�`( }�A���� ɡPЬ��k�.k6��d���f368��#$H3�0�7{�]����ݞ���Z�٦Q9���[�u��0+)N�c;�/��s9uEV�[o�ݶ��1H�J�t,���AMH��9��Ճ¾��]ϒI ��d� T�A}�Gf*-���k��kBi����������N:�f�判���*U�Vܷ0��.�t,��5Hy4�Wd÷���N?���P�����$�#LB�=3v����/b=Vd�9�s>f�(C���0Q�I� ���Q��
Je�Y�:�P�MΫ�YJ��/�ѣ{�j�+:	^C����f	HB{��C�8�M��x�/'l�T(N��D�D��l�vD:&ffEʄL����SrF�(�K��da�-�((F����EQ&�W�����d�!$t̓XŔ3Fx��V�0�v[z�Ʈ��L�	�	�|h�#ReǃH�UT۠b��@���Æ3���SX~6p�J�B�@/N/���E �H^�H
�/K���u��D���Rz�2f���LLс�yF�&fd����>�\RN�iJ����b��Y�:��� ���d9ژ�1nL]J����������g��嫭�p��(tsaWX�@��3J�U!@&G����<0L�1�"�=æ�pW��D��D�$,�fY�Y��a3�L���c�'�Iet��Ζ*#=?l	��(�ïr9�Bƚм:ϴ���Ű�aa���D�
��AsJR9B�nXJ0��%i  Q��A !!\��E�3Xʇ)$�4P;�$�&0z��f�'�qB�h��$Db=#�Px\fr ���k;5y�!�F��n:��"O��Ѹ���4,B���Tu���-�ME��ӵ4�Ȍa&��(��J�p�PfY�T�)`m�.6��T	(�VhM
�^!81Gk���`�0�����!�H��J a8F��O�H���ͤ�� o�2L7�3��եI@�h��H�K[^F�:���A0c�K�ӏ軒)�����