BZh91AY&SYpcR� )߀Px����������P8y 1��A@J�M=4����3Q�I�4���b=& �&�� �`�2��HH �'�h�MOSڠ�A�� �i�9�#� �&���0F&$!����&��Sjy��i� ���7V@>H��@e$A���!�3h^��
��2���m�xXB�hYfX@h�N�H3 j���Ύ�/������ٝA�Ze����O�/�o}�t�ۮ��K׈+�����9���#�q}�S��,�j�ɋ,J��#R��vM +4h�1�6\�� ƍ��;���G����	�z���C�����R��x���Y����*ʂ�#����Ds38�n��k}F6%��>�b�3���+SQN9ڏe��3	4�-��z������,<�j)^�n>�b��3`�u�imэmZ�,�}4�P�ދ;�w��s��\�z�KB�G���of�m��B�m�'�-B��#�
��T�K�Y[&��ԍ�.S���2�c��G��F�!m*���k�o���M����iO
����qFO�
�4��y7��Z����Bk H����>�>�&6��:�V���^=@�!7��"���:'�?�HcB0�G�BAy��ܰ�*a�t&��+ �^u��v+�uu���`��kfgƁD����|-B�!�V���A�]�I=T	Ye�)P�������B"��L��A2�.)�]b5��1Jbu������&Nu۳�m���������z2e�T�B]Xx{�Y�@0\�PɌ��$�6���Ϡ$e��P��CE�O�,�,�5�L���A�[��A]z�Ҁp���G[,��!��!׸���G�(��6�4��:���Ę`Ҝʅ���M�I!i� $q�� �����t���Xz��i�E;J
M��Z%c�C�4'��s8ŀA��D#���=י,Q q��#>����1��Be���ZI	���A�8��T&)�UZNg��9	�������g$1�k�J���KWTp(3,�`+��MC���p�-�����R�mD!!���/�I����h��[h�ͺIc��0�H��O��W��SsI�� ���44�"�r4�%�H�~PV��^'R����2�2d0hW�h��ܑN$Ը@