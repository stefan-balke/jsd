BZh91AY&SY٭\ �߀Px���������P�q��H9� Jj���OI����   ML��       �DI꞊zF��m4�@�  4�	���dɓ#	�i�F& �"�d4)����SM O�=5<�ā'�	@��"�������pAF�RI�_?"Pn�$ �hU�T��(9J��#&�v�vއ�q����ķ.:�L�|f�%>m�KFյ^0�����NdI6i�7җ4T���z;�����E�d`���H<��'�G�g'$�
[�ζ�"�ܤ	$�$*���_��sc�����DÂHi�����;��"�m��=�I]�Ά4"�Lr��+B*=���R���O'���u��ܛjҠ�Ƃ��R%���Q"4-�-&�� Cʐ ��j.��p�袠��g��^fn!K���"�.(��M�4X�1f	
�}�F�P�N3��Q3X������� �`��j��2I4���.��bB1��Z)q6jկ7�Y�B���Y��b��-f�F��tr�Q!	KRI$�@Cɸ��~b9{�NY1������YXH���$���D�⼥B��&�B&fL����*Xb@e^I	Gh�AA	h�y�_�;�L�4Y^L&\�� ��ke���5�������q�^"�ިn[�z��X*Q=��e�WR�gJH$�'4L<��0� ��ѿ_���? �_H�G� ��\v?��v�H;�A|@�����Ҽ�Ҥ|G�3�Q�0�����yET��3$����9�I;��*��$i:l�:5K ���d2ji��l7�$3�"@հ� �B��p����Y�C�rf�B��`�@��5��B��#������	�Iό�Y%�ET���
�dH���h�d����r&��G�#x2�[��eZs�1I�̱`�s/MAp�R�߷b/X0A�6��'h�:G��c0���!����f	���)焣�	���:�HP�kФlh#�;D�d*��@�xt���Xv�'�����x�� "1��x����@n��nfF�l���	�p:��Q�B��#�۱$g	�j&zhV��Ga`\*�(\^�D�xȌb*x8�C�x,5�iA�um�T�)hm���D��J.�r&�([� �fe�.�I���Y���t��S@�:"8g�R���=^�m&�� e��,h5$q$VkW�@f[��$�&6��"�a1x�0��ܪo�w$S�	���@