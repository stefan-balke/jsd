BZh91AY&SYW�� �_�Px����������P�y��p�C	MDOE<�Sj=F�CA�ɓ@hb 54�F�T        $$$�=��D��6���P�~�����3I���b�LFCC �#	&��2h��OS�&�@ �d�K$�� Q�FHJW��:4��hT�, e5�So���cIa�I4t�N�2�3}��5��۹�q��3����gF[A�Je���n��;���Q�ے�6٣�)�R��">4��������o�Ec+,3�7�H�<���ȆU9K6���*<d��� J���8�a�Z�V%���gI�N��<����f=v���,;ζ�ž��]i��ޮl�jEՑeJ�����`k�����>�}_&w9�Mq�F
4yY4�MޭF��c-xf˱_IqTwoHYM�fզXm<�7{��d*��b��M�גX]��j��&���J�j�A��+{�w�S{L<�^`�0r�C*�@M"�̨SjC���<��ț̈́`F����L�EK�N�'���oV�m���������9P���D�D�2k�uL�R��c;��2!lw��eZ�gIB���12�� ��j�s��c�Ic�����q���y���n�1VB!��EYUv�~5���,�	��#Fh����A��6�v��zd��d削
Y� Vm�_k�BS��C�b[�3�B� ��O0f�nP�I��ם�'�b�׊J~	4/P��Fv�j|(��CE�6�n6U��ŐA��RO�T��mTad ���{u���EG;�Ū�2�6��M d�`��U!J��ΪX^�������]��e\�aN���0{��L���$'�z���V3طu�Щ����#�h��M��DiR/�д~�7�-ኚ��:A�y�_�+۞�p[�� ���^=��2ߪ����ۼA��;�h�U�}�P�N�Ĭ#�
�$�"s3
Cs�oH��m���|�:$#���°��2��R���03 D�$	�~�О궈9�R���J���C��ۉ��O������3���8�d��F@4\a���A�s*A�P�گ-9�������@�6��3���7H���*τq&3^��!�8ܖG�VN�5'm�%B
H�0���/�K�	�I@�۬$X4۪Ye%D%��>摟���3V�H�p�4�Pr&XoX��H�����I���p���AxsB�Md��]��BA^�P