BZh91AY&SY�
d �_�Px���������P�t,�S@JMJx�Ƥ�Sy"z����2b  sbh0�2d��`�i���!�Jd���4  �    0&&�	�&L�&	����b �z)���@ hl��B{�"AD��A����FA�hRM"`2M|��f��x�Uaf��0��kauj^43�g�7�D_�P�ܔH���(����܉.�D��y1���Nf6�r����a�.1�F8�\�xv�E3ү\C���ix�&�l3]J +��W|�AO���( 4����.����/^��k�|��や��H��Iy�P��y"ϓ	e����ŖD�LGD��seM�>���:&��\aK���^�w�0��:�#��-��#�b0/�±R�Q���0.qL�%J��<��1!	K$�P(3o\���æ4�
�rG.F謆��
���%m&�EJ��(� �d1K��.I! ���b���&ы�dߧ�7W����ᨑ��4�<sj�ڇ`��b��T�8'1�!�CB�!MV���%}��]9e�L�[rW�H��&�c����0!H��@hN��׎�L=��A�@|W�!��|�[rKҜ� �F�l>�$2�ƈ6�$�R�f����� �-�I<�	V����5W�Z�[!%�|oj���Ț��&a�)TdxP��1C��.��2���!-%NM�p[�? 4�~���^jT�����թ0`p�q[I#���t�`]��d*��K���ٸ�����g(3\�Յ_f��� n�ԃPPZ���H�M4�/V�̳�������>�9����a����3�%�{�����s5��霣A4�� @I���B�����Ơ�"
ЛQSqs*M�P�*#�%FJ2ݧ�z⦰:�I���vd G��n��� �9���b{w�ph=��Q�,I�2h��È@��ziXE��WtT2
�4��!�p�0v��5�o�U�W ߆c}�X�BjN�![��0��!���A�� �P.�/�Ă�t�P���R4K�K�H����8�L^�~�X^��,lXF�#���|�x���ʖ��f���fA(iR���"�(HX�2?�