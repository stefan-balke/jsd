BZh91AY&SYR-�0 6_�Px���������P^wTJ�Ҵh:!)5OT�S�Oi2��SQ���4�� �&A�b�L���a4� 0FM4�"h��aF�=MmA��� &�sbh0�2d��`�i���!�H�%<L�0��~��OS&�� �42`L@��"�@A`����X��|aZ�B�I���m��B��@�Px�L����?���+�qq�������Pn���ݪagF�mE m��*���:����ߍ�y�7�8��CJkk�����h�+�â ��X�"���̡~!I�:�Y��7v���T6A
!_�۰7d��5`F��c�YW���t��\�QS�/E��2x�̐�TD��(mu�r�����<+��DR�8��ȼ5�Ǚ��
��Ir�J�i|,��$��cQ��	az��K��1C�H�BA]��,��>�2ᯗ�feL�d�J5ȣ�r;�B�)$��g7���I�ˌi�$�W�G.F�)���XV��h�1(���bB%	�JJA�����	�S	��@�l�u8�
Q�񔿾����/�[��𾹼tS^AE&�UvS��!���$�U��{w��Ҝ�/V��$Xg,�گD�b�j[�?8\����&�T
�1���L:ŉ�\�dM����^k�2�^*�}�X�ͧơQ3sr���4��j�:K�b!o\k_�s�+��L�R�Pld"��/��PL����M%�D���IN�%�g+�C���ˌ�����M'Jq��E��Z��j&��.'��>_j��)B�a%�$�5G��u����	l�y�%l�X�����ea��l?���o�Ay/ж4� #��6�#�k��v�ޓFkK�ׂwi���_0��(��#<ˉ�E�d�&��\����� $rҠ�B�nt����C ���"¤ʓD4T=ERQ6D`u�;���jB�pS��BD�#�^���bN^�Mޔ��̺�CBey� �!'���������fd<4�ˎá`����C@Pm9�g$1�aH�&8�7F�6�����d7%37-B��(���%I�0�5�C�A�bT7�����\�K#7%*���<%ܧ�ix����&��G����6
E�ɳ�g$A�|�}ͯy�R�l�h6�A1��x���"�(H)ܘ 