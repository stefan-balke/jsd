BZh91AY&SYtS�A ^_�Px����������`?y�A�8u�HI�ҏHzOS�    � Mi��=@2z�     ��b�LFCC �#	�Bb��=6�<Q��?Q ����@s F	�0M`�L$�a2m&�M���F'� h2i��v��
�d$�I��d+����sZ�2hT��Mz��m�xZI�6f� h�ڪ$`,�__�u|���#������׻c�]kW��i�o; kf!����M�y�f�Ċ��8�l��M3�
{���?��~P���}����;�6�!�vCq�'F�|�s����W�a�Vfa&0蓩<EM5m�������|�|�b i������qu�e��/��1���1�0K
�V�W1���`�L�(c��K[}家�D9�7^T3�c*x��xPm#����a���i���Q �5\J3�F��nel��-E��c)ʖ$I��l�@Wf�"KH����>sN2�	�Ca��(�6V03D($-���F0�)6�Z�鉄��(w����Pe���3s��.	����6��[eT�)6!� �u�H����l��,>!v� �	[
�rbѧ_3�61���m����;��<��B��#�
Hx��J�Ix�����B(ԩ^R��I;ݔ�U+�^eF��������5�^�PP0�r[xěm	�l�{i��랍2�i���0Y�}��7�'@8��[-s���=�@P�`>p#;<v��	�MU�W��k�BRD�TR�4�ԩ)k,���̐}�y�����q��?Z�E�c����W�ۿ^Iy�����wj���|���I�_RQ�8����S����UJ������3���X�2��� 4�g��4Q�ս��QG$�@�:v�j_"��ƇDR��(����ivv���j��3:�� �cm�� s����*�ݣa\4d�nhsK����a���͛��K��ߺ�=(�:�GV1����2�\�+�M٢e^l���s\�=�΢�;��i���b٩�&��D�V+�>��*цkߔRj��arH����v
���%u��2��u�S�#����]�E�n���P�@ Q˂�(VA�;��Ʉ��Y76*�/�_����� �jQ\6C��%n����3
b�T�]ޏ�9���>�2n���f�Ge��*'�����:��mJ(���@�f����9�/9�I��>��T��*\�<�5��kE�ɰ�z-��N~;F��ugFe��병����!��j
��0�4�2�<Ƒ��+��7ٚ�J�MH��\67ԕֳ�G%C|����	�tYѺ�oF���s���?�����N�'�.�p� 觞�