BZh91AY&SY1��_ D߀Px����������PY�l�r4h�	DS�Q� �4��� �JmP~��z@ h  d�  �Dҙ4�F Ѡ2  P�& �4d40	�10�!52i�cShR~�oMI���4 �i�� {�H�!X`����пp��
S�&K_���ne$,ƅ�ʰ�h�ԤD0Eb�۸��8M�ќ8�茂��,�9�~v���T፷ЋM�_na,�ۤ})�6��d�z�0E��&��SKeu�D.�{�0@�]�Ԡ!T4%����˳������q!1����p�A�Í΋!n�'S~͚M�qx(�MS�:���+��ې�G8a�^31J%ۭ�2��`��9��e�䙘��*��C�_w:Î�QD(�T��Z	��Ct��[\��x�J��UnF����F��J#;�:���h�$@�2F��!�m��1��qM`�d��� ���7���hbPA����7�^q(%'h�IDZ��bS�qE��cj���#%��,�vڰ�LrV$��0��-;I�6����I�}���Ep��YݐΏ\�rB�D��,Nٕj�FІmǿ{ҕ-��x�R�k���N�5���{K'0fo˚��O����zƅ�� ��i=6�{6_�TG`w&�@k���"C��zK�X��!|Q����@�Ĺ�{䪄�f��������'�`��,����in{�7���29],ڢL��34���)d)XGq�J�{J����@��J5�B�����<��F�1@P�C�;���x���ɨ��djR���=�	�Br	5�<�,�R���7�.�հ4��z�օ��ֶ�|Q�4���,�-�b԰�]y!x�: ���h�g(tO@j*�T���	���u�OY �� ���m@�
 v�H���%�,�S7���R���XAT�OY�~]A��	즴.�0���ĈH����fթ�6��b�h<�XЙ^'��$$��M^sڅ�M&L��ZT�|�C��|�����t@��$@5�1�"c�`�tfLf�����-��"��	�;n�Q
��7DK��H�
Mn(�h����\������J�1�T��1�ybmi4�܍�kA�)6�� ��7k��n����+]�1g2��_���)�����