BZh91AY&SY�jx ]_�Px���������`?y�]ب�]@�P�MF�=M� �    ���"� �    4 9�14L�2da0M4����$$��~�C4�7�hA�@`L 9�14L�2da0M4����$��=*{*{OEG�mM#M 3B~���
� Z"L!&Q"�W���sQ�0Щ0�M{@�]���hhYL�&����#1 i��޽�9t|.x"+�z����KZ�"�4��/b�!p<9�����gϤ��7ͽohg�ԧ�T.iЏ~a��o��=���ÆHd��vw�E'�zCؾ���ߦ�������dɝ�(��/I�=b��*Z��~�}�_|�B�"1S�!G0h�lh���i�J�Z`đZ,�sUu�j�4jb�\�B)|o~�M�5�,�k!��)���7p��P���:jNޝ�bӻB6u����A�V�yT<f��{]�c�EN���ȌR��TjDd������*!����±�XԣF�kF֯-�P|ab�pFX�I��] ��@ig����

�j!�R8J��� EH6G�p�W�Y�iJ^dv1y��-��.#�syc
&obi�G�v*��R�]UUUEH,�����=.�׽�Ry�T�K_$�rH�!�$��e�4�x��5��T��j��UT([PP0�x:k})@�MU�Ե�����V��ts�y���D7�����у���_S�&�{	�%�)��b`��3E0ϣ���uh���ם���6Q-���i�q���s�G���y#G���б��x�IoG^����)hl�~3����)�)'�4�OTѷ�g둊S��I_�Q.�S6��K,��j�V�`]�9h��+sDA�x8�P�".W-�SW@ˉi��v�5��"�J񳽞d83��8��"ȨJ��޳#��Ca\4�743n�%�+��'��Xn�(��)-,�i��U�(����ӟ�3�*0����o-���r�ֽ�S�鯷y��h�ݭ�ލs:E���m�ue�<�q���mI#<y ����G��2���Tg���n��w`�Cj�e"���1�E�nY ��|}*��|K��It��&��wdv��ȍS���n�;S���"Vx���w%��\�}.�d�me���Y��잉�7<�W��Q)����d�A^�QRxQ�ϊ���id��si;�O���`��|)�ڹb�*�r�����۱�L�i�,Dc�ul.'Vh�l�=m�\@`ړ }����ԩhrbq���B�,�{�6�LaE���0�>��c}IQ6��=���43�̙Ά(�tYǕ��nZ����1ѧ��塚���[�N�]��BC E��