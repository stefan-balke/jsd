BZh91AY&SY�
�% *_�Px���������`���Gm  D54��z#F� �h � ��2IC@�&�2 M4��2���&L�20�&�db``�����      0&&�	�&L�&	���� �К4�I�=���4��SS'�$�2�A �$`�� |����B&gHBE[i$�!�^'�m�)����c@4qta �"g�̎�**����"""�Qb���mh�6�S�<V�j�C��ip�&!��k��1��Y�lT��V-T͋Oڲ1��V��e��"�,$[yvd�H���p��>b&܆�����F�L�,�A�ŗNhIln�$�^��R��t�~�_uͷ���:r(��C����	,��aG��D�&EL�'$�zϢ-�960.�S�k�(FKh�M��� �$o��o���2��7�J���s9��3�'Bv$�1 1VrfJ�'&\
7�&��5�� �/)H�	�"�ֲb'�]SX�1itAKh�.BY�pP�0�hI��Yp�p�KzM��DZP�ԭ�,\�k j�C�)z���Z�X��Ky��K�x"�(�Q�U�R©�e�����X�cs�d(PE���ZE�\*z�W$R�����f��2!2�(�i
*�eF/��A����0�wNh�(��UV��9�o8�����J|�o��WJV̔��)�A�bd��aY��%��݈�S�@�b�$A�Aɲ^P�xKiAAP���ޜT $�/:ғ�2`%�\w�� )$�C�O>�͛zH03��s_|��F}:�Ǎِ�2��m�_|�8�r9�v��vT��f�&�f��� ��&�н: ����v��p}��FE�c������NGy��͈��2B ���q���]�
$�!#�z�
�Rg3A�xئCP�(�K ��glؔ@E����X0I�Ѝ'�A�ٌ��E	o��A���66t&BL���"��H�aJ���j�dDt���.*�b8�C��X�'����=�&�4�;�����|i�@0b�B�H9莿5~��Dj$#5*���c�����a3����a��tۯFsRI)���,H���W��TxV��j��3ލb�=�-�]G�i�\��ʖ�H&1ɢ$J �c��v@�� RA3��$�;ls�������T\���B��eI�%P�*�
la0@ws!<t�f��!�
����R1W�(b<������s�s�n���\��1��A��@Йf��g�E���zѼ���X�h	B�Ю,8n	��pݾ�@N9D��:f�lڤ3^��F�L6�@g+IP&�� ���(�q̙�L�څ�\H:�hD��	��)���v��<�� 2��y�ZBܐ##�J��Q�$_�G6�[D�6��9�l������0`���?��H�
!Q��