BZh91AY&SY�.K _�Px���������P��;���1�  J���dl��0�h��h0!��Sѡ����   � ����d��ѓA�h  � 0&&�	�&L�&	������&4���j��M�j���� #��+���!&d�!_����lG� �B��`�M~N\p\�$��Ю�v8��J@E�������ۭޖ�se.<�a~z�iyJ�����j6�C���>P�ms��n٣hpAC�\1��i�Qz�;��j-����Ğ�OT�!�D4G��#H�JT�F4��[���{Ѥﭵ�A~�5唄��h��Mev~�o/-t��Cb i�y����rDf�3�m��_�{�V%�aE�e�*ڿ��ż�Eƭ|Z��#���� ��"���*�6�'/�h�s*��e���)����)��tl��&��i9d��2"b$ɴ���j�U�4�ʢ&ok.��%:L�E�2�0
��B6ر�(a��$҂fҘI���"\�UA��*���q%ˑ4"�"�LqVwfU�}{S��2����]օ�VqD6b��e�./�tU)T�Vꪪ��Ae�^�Ǟm�#�B�x�:%J��-h�#m��n�5�⦤5V,���gD�T��HB��dU:aj((F��V��66��jg<�M�}3�+m2��8\_����E�ېly�V������Th���d߮�!L]��":�*1,�)���	X�En���=<�N�����G�սP>�б���Է��gzbv)h_�e�M�p�?%<��I>~Fr>>q��g'�r�Nt3��lj�!��B�C���C�Å$�8�Z��Z�y4����(n�#�i;-b�1�h;i�L��5���U��䱬�~�C�?;�kN �UJ�U*���oC'�2����_�57�R�L=���̷�T�q8����z�W�f�=��x��brr�����y��b�1~��>�r6�g߿k�{g
,[���6+�{�ǟ�Tn�RH�~p>=�B����}uG��ܺ�%�M�1ż�����p��&Ņ�w�#���VYj�lH��1ƞ
f�q]�Z���cKX�ߓ�y��ĮW��x��h�И)L>Y�nrm�s��~
~�G��*����׉��h��u��y���s|���{���5z�k�]U+(S��L��iXF*�&�td�]7%��t�4t�lnc0�}ޖP.��Z�T��6�-jdtɞ�L�=l��i�(߄���õH��^9T��Ξ�]C��3q�ˍ3c)Ϧ���S�s�g��Sz��ED׵�՗�rE8P��.K