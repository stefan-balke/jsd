BZh91AY&SY|��. �߀Px����������P��Y�4��	R������M ���� h 	M&$�Q#�4S@   � ��F��G�Ph=M�  @��b�LFCC �#	&�U?6�y3T�z&���bzO)��	�P�D�>^ox�y6 ��4*��@�k��Y��d�hX�1aѵ��#I��k#��V�[e��{�G��N2�:Ȱ�|?)m�z���ݫ�&���⒍'H@��=���YȠʋ)�U�I�k�/!��ga~�z���d�3_M� f�4Z0}�8#��P������x���4��y�z�na�u�f�Uچ�.l�v�EW.�:�\��>���[�	�Q�]�c͙�
:�I��i����И�2U	ڂ�Ti �>`5�#��䋈!U^Hh%$$��&ma� �4dp�q��֕
�%��0��f�F����W0Z`|˼��&�u�L���I�-}f	���l�u��k0�5�A�H���:��$!!�m��"��\���n�G*��NFJ�%�	saT˲�!������:Cc�#$rQ)�M#���@�H��R��aִ��lZy��7���.l1����x��%�i��wVi�&]�
<*@���_����U�x����B��Ȍb�@��?!L���E6�C��ľ��VHH@@	@@/Gc�=�]��EDI/��H���y�*q^#3ޒԉ�=I�����dQ(0"�u!If'��ɐ |��)'|�4�vM`�[��h�j,�!3�����2jɋ&���`։}�V�i+��fm�%��,0]�5$�q5͐T��X��F��ZlS�{OP}�	�� i��362K��9�GOdn<H�Έh�2B���4�Qn��#�����V[.3H8Ypd�@⼲C�JR�3I�Z�p 6�xzN�9������a����ܕ�[H���;j��(@hPk�PE�;��Ά=c�1!��#���D4Q#Y1A�.�BL����Bx�jA�oD�f��������fJ�@�24�f���s�hL���pb�@� 0@�h1�.;3H0	��傰��u�;��(\Nh�C(c,���$EǾ��ȸ��T, �X�E���TJ�%e�	�-�p f\\��(����*�VV4-�;	*�4l֧��0�z`f�`����b"Tf�(�|Qv0n�M����UW����`Э���rE8P�|��.