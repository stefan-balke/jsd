BZh91AY&SYe�X �߀Px���������P��B��C@��OS�ɧ���@    	M&� D�zA�L���@  �!!*~�=M��=&��� @0&&�	�&L�&	�����!6����P�L�� �6�2�J�,�2��w��U�h��hT�J�C)��?�$=�1���$4r5N����ݦ��[��U��6Zp>��4eZC,�S(�~���c��s���t�: ׭-|1���:��?X[$E�4p�X�d��̍(Uӂb9�3mk0��s� ���?��V�u���p����bu�T��ͫ�6���#5�N�t�nZ��nV7�	�;�%���R���*ܥ��V>�m�!���_V:4ĩ�3Q����K,B�wo9|�$&����=�6�	���Kt�`�Շd�J��/!�L/f���cb�k=`Ȉ)
�֖���ig�����{�5{Y�M��k�I�I!-k�A�����h�D�C#Vw�x�)����m��$B�{�<�/!�P�D�D���m�3�'���T�1jm����2(˲6�D���U:D-�"nL�B H1GFc�|��y���{���HH�:8�9B��.��8�2l|(xS@74	K�v��I�@�^Xj;񃺢#��|��X���`�޹#�6uq���;{�hڨ��,m9���7ss��iKC��<9���)���I���)����nn�����)ʆS��e���
��������J�&m}D��tH�Ѻ<���".W����ˋ[F��C8@&�eI��(X��X�j�0�G甹���3��)%[��ż�ǽ^����v��4��ἱ���vld	�8��6�ۊ1�f9y'�h�Խc��Tc~8����q���m���lR��6�3͖�7DG�N��P�b�s��WɎ8��q����A�ur���}"��Ǳ]�F�N�6-�I��lu�m1�U�/�Z�.4�l�("���a�!=�\�F����L�}�;&uFG���k�kϏ<y�ĭ�tDv:��Lތ�\�x]ݑ���������f��OoJ�S�Q)��wQ��񍂣QE��p��`/`��Z3���&��M:�UR��:�T�J�ʺ/V��r`����Lm�9j��Y\�~%��ӫ��F-WJX�k��eKC��Yi��,�:�]���ͥ�����#Sg�p��RR=k9yZ5�s'D��.��q�q�a�U=�3�~�ڨnQQ4�wh��rE8P�e�X