BZh91AY&SY��� 9_�Px���������`�}��q�s��t�����UG��6��zL� 2&A�@ &)� �     4�$"�j0��F�A����Jz��� 4Ɛ hM44  �B�0�щ��4    �L�h�&OT�b�Q�~�  =#OQ`��"!!+ P#!���"e��HW�f0D	��8��把�XL�I4w�)0���,��c������7tw�;�K�n�e�%���OF�5F�4�28�Z�4w���J�=ё���A��g���\�q 5�����0�F�[
���t}�2]�b�_�Ԣ ,$��?t�(0�A�1ߎy㮔�����w�7�L��$i�Z}����@�3���|M�N�ZBC��Rf�&�m�-��ڣ��Z��U�C!�=(`�������+pqR"TB�0�P���=�%�E�b��h`UA���C,�M�r�E+YRLDb5�փ6���N��o�V���S��2L�H��Lb3�b�g�IB�����W�	�"�8A����Jr!T)��� �\V� [����V!N�0�A8W,.�ybr�s�������"HP�n\tv{B�� ĉZ;�HP�UԞ�U��j�$�4*8f���vQt��%� ^��}"2��i�����N&��Ybm}24pQE�UV�	$�w��x�#�a,ԕS�jP�qsU�E�l"P�!$�(�	&�"$f��&b:IfQF���	b�1Q%�AA@��K6$1�Z��Ʃ7��G;��]l���2<9��LjQ��a�A \� ����P+�lv਴`�k翽�'W�m��$6Є������j��AK�	�%	��J�'HJ���E����B�����5�*�2HU0>�Q.�2�+����ƛ��T(&U����4�C6���� �{�O]���iݒP�sB:ݚ��Pmd"��a��$�u&�3�"`�J�Vab��[P2'��یwdXQTB��VаW�~ d}��4��j���y>��?ڻ6&=R	/a$q�9vW���L��n�+:!n~t�[�%3Q3�3�_����n�f�Ն��  #�~���Z���҆��mT��9� 4v����@���\‰�̘dĉ̸+�9�2&Z� ��ٱ@��+"���D��uf��*Qh�x�H���J�z�wo��� �&h��B9�		��ya�l�,����ؙt�;�� Y�Lt	��9BĄ!����a��rfB&P��^\r=���p�y�L(6��3��Ш�I-Bzc�a�o�V\�	-gH�:�ԝ�q(�0�A��5B����$�Ќ%i�6�l� ��*�#=�R�H�l�
�d��h^���cI��FrD< <�\���*���fe� �0hQ��u?�w$S�		�;pp