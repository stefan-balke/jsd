BZh91AY&SY��h @߀Px���������P^q*(� 2 �(TOOI���mOʏS ���4ѐ =M ���&L�20�&�db``����SyM4�hh  M sbh0�2d��`�i���!�H�@�&�aQ���  h�=OMO)�0C� �T(?��<�f)J&*�(LJi&I�#�m��Е�B�#(;�%$a��q��m[7z/��a�[q�X�H��>��e�5�8�R)JH��7$�E?�ɫ�\C{*.#��Vz3��3 ��Vse�3F��ix�f�e����-\�*H��H)����$�=�}�����2#y�m�C؃d��)�UG>����x���0�s�Oy;.Xo�$Y�C|ZR���(QE,A��vؒ�^��54�b�f2+Lܼ�(Q�)M/��R̼aa�E��Pi�<��iF/V���e��I�.���L�8ۀ��k���T�q�lcc���h@g/l����w�W&�J�W|��i�bTܲNJ?3F,bI�T;T��Lb�\��E�a��+HH j8�JQ@B��*���HM���K�bW�4��������ea�#*��^��A9�z(�Ti�倳�ɒ
M'�ĵ�	*��	Q�|TX��rV� �Xm�t��?�8���Ql�T���x�l;����J��,���e�^�K��Fvdy�(/r�k`j^V�LcP̊ϱ�A�YҒy��l�m0M�ZZOg�cPd�E	o�6�D�@9KsB��D��╅*���j��<������m�4492�г�}�h����ȸҨ(�	�� ����$����Βi�m�G��um&A��h�����e���>C3�&r/�Ǘ�3y��ŉ���V�f^���V��lֆ�VxYWbK�Y�G1_h�[���F%����90ŁTk��v��:��0I���B�+]������h���*��#�,\�$� �* �� "�6� �6!=X�%��9�2�n�R��������i3����~Ѩ3�p>��4&Sy�9�@�P���s����B�����+xT3Ӛn�2CG�����J�ˏnaV[�mቶ��MI�~�*����fY��A��m�m֒,[�KT@�;�S�i��x�m&����y�.`d����@�$A�d�����kT���"j4+�L�ܑN$.*� 