BZh91AY&SYM��� C_�Px����������P^:l�l�PJ"4Ԟ��)�&#M6�F�� h dɓ��&	�F�!�JdDh���@�h4�  i�2d�b`ɂd ф``$i���&�OA&�z��@ �y4�B�	$��������hRD�&���fۀ𘒴hV���I�!d@Z��:q��s�yT�GM��ڂ�ID����oo;�K��Nb�(IIKa��H��pe��p�η̨�F#����S���7� 7a��ڃ�w�M$
���4�H�
/��>o}qLӏ�D� ����^���)�76hF�q)�j�Ҩ��%a����z���#5����aF˽�2z浬_jnƢ)AƁ�/�����^�w%��ֽ�1�����S=Fh�)��4D���e��5J0;!E��Y��ŇE�Z�C.�T`KKF�l���Q5��-�ݚd�e�f(�h�Ym<����m}~�A���o�m�� ��f���$qp9d���ˑ���yiL���%Zg!5z�HB��p�m*q�(QR�2��	F����
J5Q��Z������Q�M�UFJ�2�Ouz�E�F؈ٕ��٠3��>(Md%�O|���z�ӱ��h�T�d�	��<̀��.��T�i�i�(�1�����s�h���� �/��<�/��IvK� �#fx�(�7�6�	+��3Ρ����q��$�J��ܪ=P�{��6�:n��PCF���.qh�wt>4o_X��36F8 p% L���! :�k`[�)'H�`F7!�:���P�*��^�H�b::+��$Eꆋ�D,�f{�-ႚ�8�5�p�.�,ە��޶�@8�^y���V��~�1`��!-��0��;@h�+�?S�tf����A��0��D�d����K\#�%$(b�T)��vɼAp�8J�阑�MN�E��X �� #�Ov��3 �:'@`���%ox9:K�bcX��B��;�n�P��Ѭä���H�3�%ia�:�A�Z���N��A�ý�Q��F<ѡA���V[CMf&�H��BjN�|J T�!�C7���P)5��i]V�H,�a��%��$�
����ʨ�?��	UD��iw	Xh7��YTc$A�8��ͯ�R�5~��ȄF
��w$S�	�)� 