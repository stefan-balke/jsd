BZh91AY&SY�hj� "߀Px���������P>4R\q��S��jz�Hz@�Fj14�2h@�Bj�@4�   �)�)��4     ����&L�20�&�db``$�d��d���Mhz���56��z! TH$�?������U�I�L$�y/��b�B��0�h�jR�i��ב��]yO���}O�:�@��0\y�p	�����=���!�;�L��dt���#fm2�,\d9�`Ar~si5�[T��l�Gh��o|��_J�w#����������<>E�L������\P&cb��b�J�*�Ɏ�A��������R]S�tDAh��@���tk��$�1A|>�����f�b�Vd^�:2s�^t3TIERKEt�!B*IbT�P�4b
�*(#u�D��i+l�T�ZD��uZ
"���61���CB��z��ޘ��NY$*�����)���,�ZE�F���QF�)bR�5�"),-�e-�	F�bd��(J4�E���#WH`߳�(UX<q�_M�MX�pK5[��.�$r�#���TC���g^�g�/c(8L�[Theg�A2����J�C��
�!�h2���ᘦ�R���&p-V�qz��e����A{A}Q�6
	���}���f����2;�v$�4	V�� ��Y�]����.:#{T(�Bg�D��LKIN�ɝ6҇;��2W��`4�s��
����A�3/9�R]���E�̘0]2�%�$����ƺ��|�"��r.D"Ӣ���n�q,�j�$� 3O��9���7��%����������xM&�VM�]�v��8����k�h<���Qq=���L2iNe�Xnz�(ȚB� ��K"�*�t��X��hM�nXs�Rh���qQ(�"0ݨ>�t'����0���"C�.Vv&�H@O\���L�ɏ��	��:�bHO��ФPR�L���7H� 9Nrq�J���6B�i�8p!���I`��x�Tf��0a�4'H�:�ԝ�3(
����Ҵ�P�q@�K_q ��.%%�"J�jr�cH������`z�:�����H��h*��"}�$�6�f�K���P�k
��jp�rE8P��hj�