BZh91AY&SY��Y� ;߀Px����������PX�3Rq�F�%�Oh���m@hz�=A�OP h��� ���   h  ���DG�dѣM��  ��& �4d40	�10� SF�&h���Oj�S�y&�� �z�F���@���%� �����i��
�
�P�5�>�m�sX�4,�d�mU�2��4>��������h�q�ZE��r��=�<^)L�n.-s($���
���>���wQ���KT �y�/PM���5�O����`�=:n��
��hkg�)$h	�L��<k��W�ˬI�}��S���Z�b�͛�ZKކ��M�.mޚ�[
�ɚ�qQ�g���<��{Vb)������#�kEt�^�M(%0{�ȔCI�&F�K�et�a�2`V	�ŰӸ�Y`e��	:L��G�&
���P���7�����B���r,�!�X�R���61����m%rX�q��g�R�%�^���1jU�2��n�U61��8��e��Z�h�Ί
�嫮@M�ŧ�����˞6��7�-�����3�W��a�ǩS_0s�R4�k��W�{�B�)�ƫ4J��N�ȡL9B"g|N-Ko�^D�!DM ��Д�k>���
�� �˥y�4��êG�J�2<�I�W��cf�Ρ���>��$�J��u1��c���Y�6�.p�m]��k[IB��0kL�"���5ԇ>~E�j��C��CѴ,���v��h1S	v�Xw�i��PK���C!u�GE�˦�Pn�s�$n�2D"��	R�TD)X= NR�RM.���3�DLr9)h�r 2��/5k\8oCB��Kô���N��Ph!����a{�b���䐖� ���$)�;�a�!�d�.�p��n`n���()4T=E�"l�տ�z�Na.�2`(�Q	0
�i�����r˘Rebs�H|�hЙn'y�$�pz �4�^vd%�M<�ZK��@q���ׅFӢg��h�q�B&=hÄfPf[��*�+pg����,N�5'v���U4ɸA�yxj�I�r��K]bAk����V@�d���R�i>/��{I��A�# ��މ7�%E���g�A�g{k�pT���ٰh7��.�p�!i��
