BZh91AY&SYH�F �߀Px����������P��7�r�@���S�����M�COS@h� �4�	Bhh�4�02`�i����)�A�
�h  4&�� �`�2��H�Dd�f��i�l��j��L�2 hSM���H}	� (�!(?���9�9��&a)�c�f���#B�3&�U�	H���O[G\���l�Y�|2���2a��D���\��m��E���P�z�t5X�Ǆ�C��\��l?l�>4^3!�sx]q#Js �``�;�D�7��t�(5.g{�����LHU3�( �'hM��+��}��_CҡEUE�eA�C�T��Pܷ�HX9�)�
��X�d��Ί,$o��%Ԩd����H��m�S�H% 8E�r.nl���r8aGPMq���+",R}p�@���Ԩaq���K��R.\K3���4P@�*Є�0���gH!���+V�!�\�J(z8�I�!P�*���b�����/DŲG�.�U�$��r[�0$H#y�m���Bv5��/'9P���D�D�Y�!�xڴ�2�m��y}]�
��F9����d�@ƅ_E��5�]���Z<o%'���k�-�=��H8<�y��댧�h�fX��j�RFsi�i�$kaw�<\�
:�9YN�j�Z�7��3`P���-�I���\}��xw��b�!��Ƶ��B��������ZJj'�fބ�!T� ��[9ϕ�3���x؅4C6�Uw��A�-�I<(�m�L[C���v�9��P�2"\n�[�.Ě[�+p�e�_^OK7ߙ���=����bP��{G��ѐs����������3�@12c&�	#}���W�	fL�&U��4,�n[�-��Mx7�4���.��6cy�A����"�>� �|խpݵZ���׸A��@h�)�>�(����E�a{9��a��7y$�� (٥A ��âB1\�pb{5�@��R��EC�X�J��_�3�)�B{e3!a�((���i~��@aq�QO��u���r17��~��hL��r:B�IdpZ���5y��h&ys-���KB�[���ZX`m;3}���s�h�Lp`#㤨ͼ��
����E����MI�Ӱ����7DK����̠tT�hv,��,V	�0���x)�i��؛ZM#��>� ��mA"�R�TD4A�Py���9�,�߃1:�A���K1'���)�@�0