BZh91AY&SY��'_ �߀Py����������P�x��j��$��OA4���M=A�   h*A 4i�@ �4 �4 ��� zj�h  @2d�L&F@��M#4i��&�&	����2Sړ�ڍ  ����4�Hky" �Ib�!X�9~#����i*b,&P� �n��#1�����N�c f��[+V��°�ʹ�k�Z�0X����U9��6���Eߛ�#Q��_d��(�1O+�$'��Ex���W=�e(�b�x;�H����J���Z[_�.({<ey�Mjhc���{(�9��K���t��MK�^�r�ab�!.!���2�ʫg������T[�Z���ަ���h�h�#�Q*����Qm�q�Y�!�Xi�Z,����a�gX�p���61���X�m��pm6wE�(F]�
N��T(��Տ��a���F����Q1-��2�:���E�KRa3
�Y쎑���<2�n�zD�(��x�ї����8r�%�ΐ��ԓ��
-�����3(�F�r�Z:KL�(��~�a�/8>�s;/BD!q���eي��!r��%�޶�+ܚ��>u���ѭ���1LC:-��D*�4C6��~�A�C���9Ф�*������B&q.&h0�e�ZgU�!�"���|"�'͕ܓ��ӉCi�P	�D�m
|�;D4>�v��ŐT(	�9��~����11uH6� ��+���)�H���0��T�F�����*>b��5���]�Tٕ��p����u/؅��@�W�ԙ+J�$�j&�,��!�]ѝ̈́�����E)�B�a9�Ōn۶*i,�s"���PX��a�.�p�]�ص�b;�1,�4P<
����g�4I=�J����&bx`�Q1�]�#),dtXB��؄�,�`X���A��L�#��$��H�b�&1vw�AR���ZP;�E��Ag*�xLm:�5��H�a7��j��h�ٻKY���Ձ�$P��*Rv��fF�T��C�A��i:]a$R�\����0�Y���,~6�F'Ҥ��
�c�H��-+	%F��E͇��'K?6bdq$��0i+�q\��rE8P���'_