BZh91AY&SY�E)� Z߀Px���������P^Zn8�(����L�j��O4S��4�B4 ɦ���&�Q� �  M  ����@�y@�  � �0L@0	�h�h`b`�$�b2#F	��D��dмJ�D����K!^>��W8S�hcQ.�"�
]S��/��'��3�&J"�ʆ��UT,�pP��7�ş^���~�a'>�gi��@��!B{gx���}�Su@a32�V�{Z�{���;��]��?�U��
D��W�ҩX�I-��V���ȭ���,K��{�D6SD����V�2���^,�
�R�m�y�W���j�\ɾ6]�
����[����}�����ۈ%l�[�%G��eH���EM!*���+p��ơ�R3�h`f#,G�
�5Z*�`Q�<YQZ�3$�*`(J^P-����
͖�b�
���=�Z�1`tAU$@x@�e�\�H�54�[��S]�{�ic-Ko:BB�I$�AC��[��*��F������q��]U�a���YL�U��CU�iI"DN��CjJ���"ц#-� @@�n9�!"�U$��ԹW��ܓ��O%�q�?�� N��V<�%U�c_��Û�#�U���5Z~��D�*���^�K�/61��Z�<`C�}��h�p#p��?�б�����󼥡���Ϟ�g�|�t���*xHZ5�k぀�-�ߔK������R�<Yv�+N��l5S5n�+K6Rт�7�T��#�S}H1���RM46��0�E7:��;g"V�h	dT�ml��{���ϴ�fk���v�����\��<�N�ѿ��c����g��6���,1��]ܙ0���{��`�)��fx�}���<���lLU�;�
�����Ri��q��=]��Q�c֮ʣf�ש�ҿ|�C[��ц3+U_�}��z��0Co.�DW��llj�Pل���әLiU}�WŪ1;��Z�ZŴsk�����!��SK�L.);�2=z\�cIp������\���Q)�C���q�eEtQ��r�k//u�\S����0J�W ��R�8��t�p���Ȋ_����!
C\�8͓��� �rʜɤ1h\�-M-�SQ©hnbs����q�J:�]��Q��r�ꑝ��[���JO�g����Cas&���5���ͺǎ���sL2����EDϥ�͇�.�p�!��SF