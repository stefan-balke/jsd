BZh91AY&SY[PS� s_�px����������`y�D8  T��z��'�d� ��   ���QFL��   2d�b`ɂd ф``
"h      �L�1�2`� 4a��4�4�aM���4G�ښ ����j\Q!&nI�EP�d@����� �B�hE�
)����n~��hZi���j��R������Ipr:|<K�mt�)q+���Z�k�ֳ�i��]ڻim�>�D �nw�X�#}�Gr�1����q8�8�5Äz�O$5�>.f��ĸ,�O���[3d�Q�4t���eO9�KxIrb�#��Az���BId��4����M�d��A0�d1�G�߷/�4H���.�!4���߄t�s�,�[�E�}ԟG��̌�U���)
ùeb�7�6'N@h~81��a�S�O�nC ����k�����/���e`s;q�0̒$༌�FD�	TS��F�p��m���a��Cֵh���Cf�����fvi�J6f�s���a�0r�:�-Ht6��XӽlgY0Le p���D����!h�Ni�;�NI#1&-FPi�f`�![��A��)�#Zl�R��bO(�l�i�Tٶ�B��3ؚ��M��)z6�(�#&U ����2A�&JB��F���۲3��P��@dj�T�q[���6� ��坑[Fɇ|I
H�ۡ�hԠ�gv��	Mi���Mz�cx$N�%���B�;�rz�Ρx�Dy*y���W,�N���q��1�2��R6H���e٧Ccc�a�t�c�]"�d4�D�"�$lY�5e@�B!y����k���P���6��ƊB}���|!͙b�`7�IxtpϬM
�uNu��A�/ �îۏ�f��`�I )�S2s����ސzw�i��e&j1I�7�9��_�>q�ZK&������ud#�}�ݨT��A x/;����y�/�Iv � ��byT*�9�#���h�H�T;����N����*�%�*�cM�-'N��������sTe���&K��e�V�ZK�y�H�mP�g�ȴ�fgX�6661�4�8bz����[�h2)��#��o�L'��bB�Ƅ��C$�D���r说5�$A��h�)�bc~F�\�z���7�3y߈]qf�.5	m�-M% ��������1Cu}! ;���; h�S��\�5P-8�r�6����L.i)��+���"�h@f 	�P"Ad6X萍%�%H�n�9F��ڝJ
Mi`	D�q�@�^�'������0�� ��y�;�~sZ���q홰�������2�N�pXI$'�ĚP���`��	�L�`�,�>G��=��e�N��x�b;h�D�zcqA��n�*�+hn�"�u�,'P���.�B��M�!�%���j&���-��Y`ķ7Ig�%*���(�إ��0�{01i0������JE�3fR�+�M�~ڶ�eK,�����0hYn2��H�
j
t�