BZh91AY&SYn� h_�Px���������P^�; n�@UF����4��@ 4i�   �T��F��� bh44 	L�ԃS�m&��a����&G��M`LM&L�LM2100	�1M���D����d 4ڞ��R�I!�H��U	@@���q4��pDD�����#��
Ȍ `��Q26���'ſ�����:ys]�Q�x[w6n�D��������\9"xUR!֮�-j�	����y�wV�RF�p����-��	��]IV���'��h씄
�P72��K��~��x��y���t,X�#7M!�%GYDaH@��t��&E�_�sm�A�C��
�\��+Rf��i�$��<y�����N���DR�+)#YYFP]l�UsU��[��/�j�i/YV:֛
��u�P�-H�[s�9v�l�80jb�lP�qr���%��x</�iɝ�Kpl�ͱTZKc��HB[$�Jg7)����b9��9$+?�G.F�BF��0b���w���#�R�)'#ldG*��T��!a���	�&�k��o��)�,���$���O��:g��5`=�hA�	��fX}?j+M���v�U�.�Q��'�2��DR�3���p����v�g@�0�q�����) d_>���eξ�+�KӲ�m�� �F,�y�&&m`k^QUBd�ɇ���<J�I;��,����[�P2d2;�CsS&-�9B�"@հ� �Bs9��iD"3�ya���A&4�8q
����X� �v��T�q�.�?�u�0b��DWQrQ;��e�"TCD�$,�6[	��z��H�[�&���Y���+&���Z<iJp۱U�$�Sh�Á�G)N��6L-9��	}M°`L�`Ҕ�!�J�z��* .0I��A!C��llj#�!� �h<�aB0+Q���EC�P	1����hOf��G(H^{oH���/}����^���ݙ�Af�N��d4&S��9B�R̅���f�!H��XT�8�t�4��ӵ99Dc&���K�Ӷ���� �Z���%IP$��[�����P 0�iZB� �L8�WE�B��I���D1z���a���li0>}�A���Q*kV�K��L�@<wM��m[
Y��g��
����ܑN$ۼG�