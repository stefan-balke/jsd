BZh91AY&SYI��� ߀Py���������P>�j4h��G���6�i�`�#&FF���L�1�2`� 4a�$�j����F�I�4�����3H�L�1�2`� 4a�C&���6�y�Sd� ���\M ��"D��$@���AȽ/�(LXhP�d����m��(B�жcM�I��YR�g���G[��2�~Y${=��Ëㅧ�Ю5R6�����x�-��Ǣٕa#X�HӠ�Jw�3%�VR�yP�u;D`�z޹�e���@��I�ğԒ������aa�	�|��G@}�(F�E�.4���b1VBdۉ]��R��{�_(%��Q�T4��(|\�r4N׮ٜ�5�����C��P`
�IY���6�cE�pkf{�jwˠ�M���[&�֞���`ȼ��o&ݮ�裄3��\k�k>��61����m�4( ����_|��iIBx�(��,�3�G���{C�*�C"a�L�m���H˘J��$��k���b�a�=��������:������?� b}~����E��#�)H~ 5���ϔ��UZ�ԮZ����n-�9O�s\���S$�����K���y�#c�`���m�H�bi($����;���|FY�K��K����ʁA>��K�jS�2�qP���=�i'�U��4R��X��\ƢƠ���'���5be��0��Pw�P5�/�{º��gè��hgcM��cI���ahY�?`ۧ �-6)���G���M�������#}Q��_ ���1�9����]|�P!K�1���ܢY^�C�k��T��VM(�yd��k_V{P�z��������W��-�4'Paya,�Q���^Ҝ́XnxOQ9k(�� 	6( �x�DACK�"KH��L�l8*c(T�&� �,�� "��j��W\�ʀ2�~��G�yϲ���5�� ��Gr����F��q>cpXIA�/CC�0���
���o�h,:�E��V�\Nh�p�e,"H��H�tFeFc�w������fvH��BjOF��T�""���jt�[��Ae�II_
�k~�?KH���^d�`z�8�������Xb��%��c[s����mT�G�����!�BQ��A��ܑN$d�5�