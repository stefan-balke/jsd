BZh91AY&SY �֘ �߀Px���������P��pC.$k�%	꟤�zy)�=C S�  �@��L�E        			i�Q�S�S(���FA�b40`��`ѐ��&��RPL�Sz��=S�F
i�� jh�K�+�"Y"Ȍd��+�����؃
�@X�k��f�=vF��fL"M�EM��������}���R�:>�����f����T�'���p��aG�`�#�-Cm����i�Q6/nW8�����X�̋�nvd7'���[���7����#U���DI�V��H���U3�T�54��V=��j�%������ud�b�%r6�%H��C#�%��o4���?P�&�߳F����>���&nL�Gn��$Ƭ���B�r T9���֤X�*��Ed
����VdQ��Ai`+F!�fY|9�5Ȩ&̬���RZ�ʨ���(�d($�g�YX�tH�7-A)v���&J�A�o/��XQ�,�:DV/����lc{�m���BO�����Iw�ʅw�%�Z�]���x�a��Hܑ��̋��Pă��\e��J�E�}�V!�!�ny�;Us��Mp��s�xH=^�ǔaH��l�����3:p����O��S�������k �H֫:&y�͍�A��b!hs��ܻ���'�<�4zTG�Yg���\�\�y�)d5Z>Ǎ�%1�$��L�#�2���yzSu4﵊�E,�k�w��,|��+Uⱌ�j������ϋyEq�+�9ͫ�e�͋Ěα���2�l��3�Z!��Z枵��*�*��1��R����i�yZK����o����唢���l�[|#=f��.X���ۢg]��_6��j�(��-�0��T-}	DaL�	Ūl0�ݶJ�S]@��v��qQ��Ү��;�g`p�Ȯh005,�E�qF���5,��
:qPE�;�X���#�K�\6�a��d;X0Y��0$K2B�-�I�z�D���9���%�=yI-R<m��OvL�e����kk�}	��j�NED������5"���;6��r.xe4�t:�G���U*�S~�-R��a��4�9����X��a�io9�FE*V�Eg�?	pF�$:����Aȹ�{F�LqR=��d�k��weH��[u6T�N��CM�ks��F��[wX|wcU;�e����%C5O�E����)����