BZh91AY&SY-�� %_�Px���������Pr'�P$ �I�S�~�M#�h�z� ��%L�5S��@4     ��"&�= <h�  �2 sbh0�2d��`�i���!�H�$�LiOSLҚy��=5=OI��℈H�"���Fqp��
CB�&I� �M��1 Ь���)����d3��[t�:��쭩~�`�uRQ<�o��[���1ân��nL*%�������6g�ٖbf��lf�A�=��g ��'=��ڜ�iZ�w�����s*��k�P3��4Ҿ�����L�a��>�FE�!:���c��{�,sj���}��~�6p�̚񬲤"��#@�����,���I$�i�+1I�X���I�q$;�1�;(Ό$�*�&�Tȡ2�l�NoH�!XT5\������&1%�Z0�͖l��1DQ%U``�$�r��ᨍ�If���~���f���#2��T���p0.�Zb1L �$�z��Q%�E��CĂ0
F�w*U����w!4�O�����yuXy��7�?,p⅀ӛ��C�g��i�ũ*�c���(��cu�gX���ș_x[~ε����+�'���P<�\�0�(�
d2hx��श����ڬ#��5���y�*&n`YyH��C!��(��A�[�I�J���5c���.��
�.9c{T(oaК@�&e�V�G��M����.%ƕ����L���p[��@�9v�Yq�LP%�w��ƚ�L.�1%�I.����{��7 ©*�	Z�#R!Jq9F����Uv����TD��H�#��<A��9���j
�)R�%n���GI^���P2�B�%�b��$�CJs5a��9F�i1 @H�@��+"�_�(�� w�7�t�bh��yQ(�"3�Ի�B|����S��	������8@;�۰~���>��4&S�����!>p4!��1�:;6�()�����Y�.��P�Nh�x�h��Hq�Y��%Fa��"�C�A��X�Bk��e��T��P@�04-�jn �o�vK��\JKD* a���S��4��&Ɠ� ��F0�X�YJ�|��`?�s6�f�K]���`0hY3��S�rE8P�-��