BZh91AY&SY�G �߀Px���������P��v�"g�v(���)�S���`40&�L$Bi��F�&��444z��F��A��H!Sć���FP4Pd��4 �	���dɓ#	�i�F& � �$M ��&#Sd���A� 4�O)�|�\�D��$e�d+��~*����-�H�$2Z����p�7���(9L��l1[x��6�캡kgٵ�*� ��(�������B[�D�K>L�I!D��G�ZxC���а��3	��#�"�<�M�G�^f�zN��� ���ީ$+al�H��DG�K&ߏ�\{Q(@��O>���pcpdF�N�Z��(���p�2,�X���M,J�2�*�q�����P�a�����Wp��m@��ʄ�f m�6��%�H�\>���`�mv�Y�pnf��N!mHy����n�FF�R�×���_�Bc�S�L�L�k;�0���������vli��x�El����9�ޥŧ[`N4��P�[Ӭ��3U�8�7�!	K:I$�Q1���_|<s�`ӖL@��29r7JlH�(���mc��Cc�ڃ-���d�},���| ��$��k_:�bЊ�9~�%%^��8q��[���.�>��7(�����Ϙ7j�FV��҃���>�@�)>K�Uf�R�u]T���{��͏\���y��g��?�{��f�RG�Z9.��w�t��yKC��<����?�2�x�C>��ƛ�,�D�
���%-M����K,�2����7yۂ�'�H�>�r�-A�2�z��a!�A��3�EPjqp���gz��ǭ��g�E���"��CF�1�Үᔮ�����ƶ�^���ٲQIk��b���<�Xz�׶�dY�����䉺�[�2N$��^�)��_����Ϳf�����%��<v��a��|Tj��Aˇ�os�,;�6�48:͘�.�&
��tK�l��h��a(� $��P"B�.(664���*�(�FC0jIqB�OZ�Q\1���U�T��c����^�B慑��9�kif,:|,�ܚ�����OC�ʺH�0�Q�R�]��1/�{����|��J\��`k0UJ�
s�r��h�V�M\m��M�9��/AѤ	љ2U�){뉁"�H�!��MF�KC�c�}��*G[%�e�!E�F˴��'mH�ʶb�RTOrή��=�.eo�e�gk�j���2e��SR�ܢ�h��ϓ�rE8P��G