BZh91AY&SYv��T �߀Py����������`~}���y�p:�RF���
zO�#@��i�&a4S�@)T���M     dɦ�L����0Fh� ="T         "�ѦOP�C@ �4� �A��DA5&ɉ�j~���4d�F� m&�	�X�I)@�V	F�&,���C"� FuF	��0O3��]�h�52"" ��x{ݞ�g��ޗ��=����Zw[v�պ�wu1mm�ө�:�Q7��~0i�aW� u���$�:�{�)���0�m���I
��HqIc�)�t{����e�k��.T�t}Y�I�y'Y����L�8��+:;�a�<�6/�� �a�j �R�I�ҡ�p��2�$�Dm��R��e����l�?��HLm�<�>��=,<�s[���.��������[R���ך�U}����_jV��.��I2C�;�������Åʊ�o؆<"�sS 8{� |G�k�"yl2M���aȍY�M��RPp�˽���&ʋ��J�0�Z,қ�Q ��x���h�pCbG#�)I�ǌB��Ha&`��Fb���,��8.�_�&�q� �9�zA���"(�a�)�fVw��`����:�1�2L�i��h�\K. ;0z��b���@�j�-��.��dӖ06��j;"� l���b�Ђ�t�e��<B.u���G�c+ѳ���(^43ۋw,�P|�z�t��!�B����4.��Q8�U�@�!Ր�%Dcܺ�"�3bDdB�wǾ<�H �A8  BQ5�emt��F��c��!"�fS�)�� � �)DE\TM0@��p�e�T�&\�uI�1��	��"ZdXt��UIF��B`1�()��	�#7��6	6��	ȭ�>�9�7H�J�4N�����g��;���Kt1��})7�@����:�J!�g��级��Ӛ�L&�gv��ΔF�	1+��JHE���5k�[���ΰ���!Q�BAHX.���Vm��!�H.;
ն� �*���k5�NuGf�Q�@P�p`n^렢`�f��`�z�d��P�[z �Lco�t�?�v���DT���T�����4	��!�YEm
l��g�١���sZ�ʐ@�m���$�hUr�����`>�v�A�cEQHX�)�?�])��i!vvT��Q|d�����[��B�T4g+A��P�)����c +��K1H$�"\�DAq�R���G���}��o�C	�l��zH^�!�Ga^c��bx����< ,05�LJ��l�đ 2P��P"B����AC~$U"��M��^�EK�X<��%d@K,��u�F3��Tv!g%��>�^&�jԈ�/�M��w	u$tq��ChЙ~��u��,���F`��'RHW
$>,K��3 ����Aa�ꁜx�@0]�4șEGc����\f���+B-�q�K3��K�r�*���p8�CQ�3�N��%p.pYg�!{� �n�\k�d����P�$��f܅)�R[��K�;M��A� ���3"����8n�C��k�ޫ�~��h:F-F���)�����