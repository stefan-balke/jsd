BZh91AY&SYx��B �_�Px����������P��]���:4� ��)�CF�Q��� 4 $�)��?Ji�� 4ѐ@��I���0  i�   ��0L@0	�h�h`b`�$�#	�6��I����i���L�μ���,D`�2 ����j��A���+&)",���6�=2�d"����l�,l.�\�G>��^�f��w��2�h�4�,Gw_�K��;��4�mE�%)�o�Х��>�g��3�����+!0�NǸ`�Y�5�����G��R��"Y�{uBB�e�.㬄���֘c�:`��x��DY�n��\��JۛQ�M��-�V(��S^�ۚR,*�}�a�+��pT�	���ntħP�#43	2Z�hfXC4k!`����m����^�R8��cNh�4B��gx�r�����7hzWwT�b����;�*��J����K��m�:���S�S���"5��#w�ڭ����&�F�^�ɒ�G?�S�~[N��s\b*s�X⵬��΃c�6�I@��3��$p_rɀU<9r7J�uK�C�T$D��9N��T1(���&e"F7)���"5�AE%��!��$���B12��BD	�±%/�g�r��s�}FN@���Sç��T�R�a�	��lO�����S�Y�w����`R��2eE���1S��7.X�>�:D��]ή�w����w�7�RG�Z5�ݵ��ۣa�LM�-�xh���O����;S	=RG�5�s��0ؤfbc�	Dh�?+Lc=˛1��-{�^�q��A�{�G��d"(�n���titL�{B5��µ��h��!�O����f�H�(�Ի���i���W�5�ӛ�����%�Ww=G�ۇ=���I�`���(�޺<Y#�Ɏ�o�p���x�D�]��H�N�$)����E���:阱y�(�
�\��q�\�㎮↙�$::d��3�Tuv+竬l���id[��CJ�E"���mU~��B�2����d\^��;1q�A���똁�2��
���HK_KX�}���^����#��/�ВޕZG�����o;|�^�6�N����oWa�Q)�'��2.�cT*9�qX����$s�B�����^V�t�׉�A��V�*\�'}[]��L5tۋ6���W�_A�b�1c�%Y�}�$����q|�r�Vk�(:\ΰX1���n�ϝ�0�Z���K�jF�
߭���Z�F�5Ct.dn��Q�賆��ꧽ�0ɓ/�Mj���C/�.�p� �=܄