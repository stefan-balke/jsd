BZh91AY&SYѲ�� �߀Px���������P~:.˄A@	BE��4�4h��&&�4�4�1	H` F  	�� 4��"OH z�@  s F	�0M`�L$H��4&�F�2  #S&�'�HP$���`�����ļ�Z���5��6�3H��d�0�h�jRQh����:y�臗K�TY��We�!�����8�p"�v���E��,��Y��I��B^wA�ɾn��h�EL �q��i��Jxɐa�٘�;�iY�޹��8h�`�#�dB�k1����Y�H@� �M� �@�+�E�jyd}6��݁gt�*.�x�L�"�o5�� ��`��ځj���P$]�"�!�!VB����H�@"aQU5a5��a7pD8���h�ܛtU�����"�ߣz8BC�AD����*Rm�
�)Vgv��"D��aXj��,4[R��a��`�]�YE� s�I7�+����>�����7�m���6�Ʀ��"�)����	����uH�	�$JH��*`3L�%��'jM#��.�A;IH$!��Ԋ
�����[Uו��k��+�1{D3y��%� ���#�=�f>? �8Cu�5���4z��^�M�Y���`o�&p���h���v���������>�$ˀ�	T��5�t�|�J�K�2�_�^�#�ٴ�RcD�W���fð�{�L�EO�[h�@�-ge��f���E	r�85D�@\鋋 ��D��╅*�����!��.E�Uޔ�Cq�Eϰ,��@�֜-%H�`�uF�����������Ij�����F���[*��K�Qk�m�Un�#���!�K���#�d�+XI��k��:u��̆�������0%{G��l�^r�,Kx�02&�'3PV�s�dL`�	��L�ұ2 �!��D��*�p�s$Th����U$D���ݘX���=����������5#�X2�LH&)(K��SB�ѡ2��Ӡ,HH} d�G c=��Fa4�q�\X�=��]HLm;�3��ɢ�$LqzXn�Fl�ါ������i'P����%��Ȃ�Y���4�B�C���H-a��u��k[�d5�UO��e�z�9�M�����.`mJE���e$A���^F�Kh����F
�OM���ܑN$4l�? 