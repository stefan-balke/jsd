BZh91AY&SY{G� _�Px����������Pw1�8�A-�(��{T�mI���щ�=4�2�����Di�A�h      ���j~���4i��  � �0L@0	�h�h`ba"��2M�����i�~��<��h $��R�I'ʐ�!"h�D���&��pAF�HC ��xI�yHhЬeXATL��6]�����ٳ�ueH����G�G���m�n 4�#0DF�0G��&�� ��N-f!��Աa!�'B֠�um|�ʇ҃J��vHEm�d� U �sd{||%�N�ڮ`Ǻ�8c�Ղ�dU�6D�6�u,�ؼ֯e���e�i.�Ld�ޚ;�ICV^$LLJ��Qj�ƪHf�L��eq�|��˼<aR.��J��Qe��+����R��T���A̶�1E�Ɲ�Z�y�3ȴp�Q!	Kq$�P(���GG�7�N1�,������Bi��HA�ta$;�`�I��*dPG�����y��@�l�{�TEQ&ֵ��������>XM����4wA�e=�:� �A;�F���*�/��+X�j��GYi�M]��bqO摂��ĉ��w�����xY��� ��^u>ÿ-�0���oD��^c2�%/�1w���2<�I�X�mT��f�ҁ�Ő yu$�Җ[Z#��j.(�l�!3���jhd����@��n;]������@���	�H��@�1'�XT)�?�� �Xb�(������2�@�o|̘�.�(�Tp�Xe�M�HY>���[CJ��$o]� ��W��^�� ����R�vd�-L��5l��| h�O�>�����4�����ŃDEQ�iV�-	��llކA!C�B���=��Bn��v%U�1E���T$�v!�r�W �i�$���3�lÉ�	����SKG �5�s�6	��u�@T�C�B�����#�aS��,�L,�N���2#�� �q��ee��EH"��wu�RT	(�n�&"�� @���@^5E�Ɇ�YmH�j4t78�`�*���O�H�������iw�3�X���qAaRH����:6�F�:��ᘍ��B�AfB�H�
h�� 