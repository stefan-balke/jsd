BZh91AY&SYQ�m� _�Py���������P8x��@T%MB`����d��`j~��4dƐ�&L��L �0L�0�DM#T��hdm� Ѡ�C��2b10d�2 h�00	�4)���2 �4�0N�d�;��H��H���t�O�X��ơ�6
�!A-~Oèn�d ���S*�H2�=��OsN�������ΣV�"��,�9ͮjZ[�Xz0��c�@�3���>ۻfi�)��GGl/$`���A��)I�l��Α����BH���BB�>�_71���}R$H�|+w��MW�m��{;����]��wᵦ�Q
5���C��*�[̬�%���J�� �4�d����ざ8���u�LY�<�⑕����L.f�IѢ)
҉��1��e����McW�YZF��\�ϰ�61���cm���]���)p��M��C�p���,Q.j�12dT�%M�H�%��ɂd�țK}��3� �D�$C]ޣ-  ��>��Q�R��K��:�3���QYb��_��R�5��5$��D=������@�rI1��tu����D��uN/�!BŖ�7��[�X�:���r�P�?z!���Xl��x!�A�@x��teҾC-��z*+9�#L)��-�G�s^뀠���Dz�2<Kw =�J���V�z�hPmd"����-Q�nL74���V�w���t݊�>�楝��6�lN5�:6�����A��7��R��9X�Z�c���mz�#�C!A�!w�G����R3i�L�mQB�1-�1��yU�QL�L���ǟhg��l�Xx�$sO�g>cy�^�����&�� �x�w�Tz���l�^t��K��ы�j
�s���8�Q!g 	��z�,@�x�D��"�P^�U��cs�Rh����T(�"0ߨ��yS`�Wi�PC4y�D�#�:�]�ၤ�hD����bw�`k�='a�$�����WJ h�r�"��(P��W�γ��ś���Pm9�g$�.��(8ΌxGQ�w��*�+xq��q���MI濘�����jd�b��P,G�`�33g���!�x��*@�ZV��)�`��փ��irt����,d�*-2D8�{�6�M���\�5�#d`Ħ�u�rE8P�Q�m�