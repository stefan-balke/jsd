BZh91AY&SY��S� `߀Px���������P��#�8pkM 0��M=Szj�M�z�(�� d ��5=M0�@       BH	�h�ш=OP  b s F	�0M`�L$H�d&4Sh�=M?T�4i� @�j�u4�� �TP�?��1��#�^1�*LJ�&S_��A8��d%�İ�DCK��tH��=|{O94[�����o�jϧ$a�*e���\� ���d'[�ۜ�����b��A�Z���#�F�,5b��M2Ѡ��2.�x圉�0�ƴ,�$iZ��Y�By�ZS*�ơ����hA;{����M41����z�2Fl��SUE����vE��S�:����E��c��7�:�&��ˠ�X.x�6��j�(f��0$��Jj�
2�!���{��!��#P^�9Vr�<�!�r|7
D$2����PdBY�j.��P ���AD�\�k@��KJ��f|�l�
/&VPZ�����6l��m%s��.Txi.}Z
}�U���<%�J�Ic]}�䃰�s����%E���
,�Z�jH��B�j��f�eT�F0)�+g�cbJ�b���&�p�c��nmӣZ%EǎHy{<��>bU~W��eG7l���@`!b��/N��N��<�0lR��|-RIt��)Ʊ�;r��1�#���y��'���Id��)���S^��KC� ��y4�g�K�E%#�`�L��2���!�Ƣ���dy� <(�V��īk3R���لY�.�(-NZhE��0j��,ԭYȭ�p3�̱�]�C���v��-�~(1���mj�֬*<Iм���˷��%�A�)r�-�ѧ=���fD�[*&�H����fҋj4��
f�k�8�-�?9�0"%n(�&�P�,P��y����
������%���@��W��8��@���P�U4�	�KA9����3�`��[���$X,w_,HHF����\�U��Xd�P�DI�A� �� "�sv+��'��Ļ�*i��`�!�zK����Y�F�H���H�o;;�bf�����2��g ��I��`���]~��X��X(}X���G��Z.G!^vв(T�e�� ��CE�1��g���͛r�*�+xFW�&V�Bu	�;��%R��kb�Ҵ���A��o�����-a��t�����R�x���,=<שn`1$�����cl�yT�֦�,�@O��gh^FJ�P�Y���&�\��ܑN$)�T�