BZh91AY&SYqM�� �_�Px���������P�73[�p %ORQ�)�LL��4h�F� h ��)4 �zh  �F h %S��"z�i�M Ѵ&� bd���a2dɑ��4�# C � D�Bm��bM �zM�-�IF�	@���+�����F"�`EX�D�
h$��|�ہyM$�
�,����D -�;��n]<�r�s�c�ֈ�k��1`�k�7���d��7�b���xl
��LBIƚ���ҚQaa)�Y���x<�ן$���d)�[1�YFcvEKe⭗r����J�xM ��� �O��KO�~�\P&�1�_I�t�ɝ�n�W;r���h�i*)d�BN��� ��)O�"�[�]hg����f���0ft�����Sig)t�R���t�#-\����+�BѢ���^�L>F�%e�L���PvZ�fy�cXb��.����T��)��Ԓ�w�DZ�	� �D���(��E%�衯4*�#���z����|�w���R�BE,���eV]B�{��$!'��I�1�L[�h-A���^:"����$��Sr�BI"�	D$f�ʐ:).�/�e
"%]�6$D&�uڑA�� ���Wy� �$1 z7��ա��vB(oGwu��GN`��ラy/Za�a �@b��%�}:+)>v'�(LѢ0i������EJ뗋8��&���n�?]�G�
.�H�������?���J.�� ����2�!k(��A�H<��8`e�A�oIy����F�q'��LL��Y_��Q1�d2���l�qo\ؔ@E)k-%K0�:�rР��E	q��A@e\ɇ+H �0k4R��*��3`��ϧ�3Gp�m���%�9�ar-�O��{sj׼Ԩ)�O����Ƙ��2$�	#���鯈]��dU�в~�{J-��M}��PD��r�3��FN�4����3��m�`��-��r܁{{�P�Yc���@�`�.���H�P����if�4NQy0y�-0�ͥ@��¤�q|�" ����$P/
���$9��b��E���B�la����B{vl@���G�æE��	���ӻ�H�\�6x���/�����Be���б-����h�b��ځj	��3R�X������P�O��d�4I�$<
����TfYo�+B+�7�`3}�X�BjN��
 Ui �;u��!�jdN�¥��H-a�YIh��j���#��h��M�&'���ħ ^�k�֜�a$o��<[_2��m���CA�0L��dw���)��m�