BZh91AY&SY��� �߀Px���������P�uP`@��&�O(�#���@ �	���dɓ#	�i�F& �)�&�&��0�  @0&&�	�&L�&	����&�jf���L)�O)� i�y5=O)q$�ڐ�!"h�D����&H �@�!�k�-�0<��hV&U���� .�d����ԟ������p��H�w>s\Ek��f��Dc��K<�!�I��ǯ�c��,#Mb�o<�g#\ɺ;����r�)��`�t�$�L�@)�%s���7x�R���������6dFɞZ�F�,Y*:6E�byJ�:��̝�)D������ ��d�T)���+�
Eɪ+5qDpy8�0�eB	PP��$�{T�3��`a�M�1��{�Mj�324��5-T��3��c�$!!	jI$�
 c;�&�l<��rɁY��r�n�b�%��%$;�©�m!h�$(#�CA���$$5z#n@�d��C1>�,N7�8����Ȇ y�6�O4̀��*iBl����#c�t��S��X�!d�n� �t1���ΘFD>��v=+����u��#�A ���4ݤRp2/�+��jؿѝe�Jֿ�����	��01^u���D�w�2"]I'|�4�l���ѨYL�5����Ɇ�œB��D��ПqX�UBL��p��T�[�1���5�PT)�>�4��C���HP	��>���	��� Ē�"��Gj|�v� ��'!k5ó\����#������B�B�p�je�KU�3
R����^�F��#�����Nq��S���!�&0/$إ# �������$���B�+aB���~D&�0�#Fd2���D(�BL`�`}y!=\�Ds�I ��}�"1��|�5�� 7�����<�ͽ��4&W��7H�>V�p��#@I�=pV�N���4�ˋi܁���UzQ!ލᴘ�8�T�)hl�.06��U	(��o&"��L�d^����a�j��D+Q��8�ha;�z�F�g�A�I���7q5�(�$XkWDm��ݝ�}�u��g �14+s��O�rE8P����