BZh91AY&SY�{�� _�Px����������P8y��ѣAF�56��FQ�4=CM2h4 4� � �`�2��HHI��b 4    � �`�2��H�Bde3$�E<���=�<� �=G��Y$�HDBE�HD?���:7?q�!��2���[6��f4,�d�����JT������upb:�1[)�O�7�p�Y���*�e:cn�o����l�|C�L�Q��;���-O2��b`����������$�0�m( V9q��J�p+Z}B;?����˝ɼ �����+�3(rr�t�Iw��l�"s+0�DV�$��f��*�_b�[��ޛ%>�{vّ�x�X{��1��v���65;mZ�h��4�e�n���f0閲�"�QR�/<(�00�v!rh�6i���ټ�����w�܇���wKߏ��lcc�m��D!ܱ�����G*�yܢT�K�1A����66���#c	P���l��T腲��@���Ɔū��&�>���l���r���W��ߨ��h����L"}���YP��7�焷�5�\G)r��D����Z�vV��"!a��R� �T��j 0����:0MH���� �׮�}K�f|_��FY`ƃ�D����t
$��^��j�zT<{�E��'�U��P����s�5�B"���WC..�a�B�p`֒���O:kz��,5��"48X�/8�B��� bM[�������%��O�=ߵr�J��ꡣ5�G��_�3�H�:#DB0��^��djfa$�����:{ҔlG*P�\9�>��0U�vi��,i6�<9�4q)��m�5��(05��3�7=�x@��8�Bb�!�V����E�0�������\Rh�{�D�~���!=���p&5��2CH��T��<v��b���gq�dp�!�cBez�i�,$���`4t�:[�dD�L���a�.	
޺��FӢtp!���"c��7��3ӆ�b#�Mr�"�*y�\F(�$9�x�
X^Is�MW�H,�h�����X�X��#/.M#/W�#F�K���Yh\�h�-EE�H�dp� ��`���,��ə"���LE�.�p�!l�x