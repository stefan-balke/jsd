BZh91AY&SY�"$ _߀Px����������`?y�Z A�1AT�
mOSOSO(�   �  jzh�4� =C��   9�#� �&���0F&P�4Q�{)"Pz#@24��i�� �`�2��*I	��S�M5=L�I�4�L�M14�HW:��&$�!^�櫚��
� � e5�;�ۂ�I!�0�M�S�@R����߷�ǻ����C-��mkKGZ�T�U�a"o��[��<&��H�WgLmѶ۲9r)�L^�#ݜn�����m:�fS���hι�Wkk[k5�e�v7�C\�Z�M�X�_x�1�b��K��g�=�+j�g��w�uW�%ր�L��� q;j��z��B�sHm���b.�5{���:/K�k=�V�]���}6���O�:��]d�F8�ˑ�a�j�fI����f�t_;��OY�"�,��p�R�~v�LK:���k� <�a����h�fek���a9L�fA�f.s,00��z��l$�2�F%j�X�����,��Sc����"6���4�
!ڀ��S�@�@�w��dM���"A�$����$�C��ʚ���i�	4(hEƦ6),� �Q���Kj<���k��o���m����;l|>P�B����B��m�Z�j4�&ATU��������<�.8F��H�
$"�m:�^VXj0��!l蠠a�.-��ZxqO��O>q0��X`�,� B�����J�
혷����#�f�����<v�:@����d+G
c��9A(4}��V(��d���ht�흾��oa�NN�@��B��K�]�^Z��)KB���=2/ˮ|˚I�=>1��>HΆ:��d���s߀�},�<�ROk�c�ˆ&��G1�טy5vDK�Z����ˠ��7�!2�B5��"��gǎ$83��Ůg��h���U��t�13y�6˟$��m���v��ۆ�����T���]�_�7ys.e�2���.�Wa�yxqa8�%�ҽ�SG�_O��-��@��<Kb�-��o4�v8��˞)5MxY$n����,;㫬o���ح�&
ך���r�#v�ό�� �GUPX��V���t���XgA����\Tс�c �]�(�;��q�Yx/o��:!f͍aeH�����K��3Eë볃���G}��7�%3x���8��6¢�K(�S���	�[�v.Ǎ��kN�����ʩZaN�u��5[u����7o���ːX�Ɓ�T2�"�*zk�]f�������iT�]S����š��y�#����Q�7�M��~Ƒ��|ܧ
��z�su���$\��hf&ˢ�l�z���Os��y?jmu��TM:���w$S�		��"@