BZh91AY&SY)�v� �_�Px���������P�r �F�!)5&&��~���z��Ѡڍ h ���&L�20�&�db``� !S&����L���h��`jz�!�	���dɓ#	�i�F& �"@�&�	�S�z���'�� 0S�^My!
Q!I(>���r4%�*Ф�%0C$�x|�ۀ혀�4+@��p��Q*A���V�c�!�ޫ���߇4�[l흁ciD����n��Z�����(oV�iƤ;[�=}���
]�e�X�j�E��\���*=$��h�WlH����s��*ݢd�P���kE�?��(�B�Y���ã��1��B;4�2��ݺ$v����1WHg,���[�W��u�i��Ƣ#�A4�li ���̪Ư�j��)1p��A�J�ox�� +gdP萁�#^� R����1̂P���,��4�k��oz-*�X���)%cK����|��qG��G����A1�+Sg�U�tl%�8�t�,��B��$��A�~'�i���4����9r7J�i+��� �cD�E[I������R������
("��3�&$$5�W"��"�U����ߣ�Ÿ���]�!"(��q㪊��-g�;�xs�����pt�6n��l�3r�62V�E㕸��:�;Kj[�?��M����TA1��5߬S�d �@}��l�[zK˪�}��$jf�Ƅ�S`���|���P=�l��޴�*�٩��f����Gf���E	r�2j�2�ɇ�08��5tR��U�s��p3��c��P!�>$�=�?0H-�
����B���d��6�J`���-䑅Q�z��3l�!l�)-��#�s�"J��	�BX&�v:�ف�NTq�������h^<~E�og�iiZ�@m�@������^���h�Ib\Q���X� e(b��r�$�2� $zq�A!A��t�b
�Bl���s*M�P�J�6D_�R�ބ�SX#��0=���y��`�`s ��i��R@b4&S���!�h�0g�`F��S:,U�c���9ś�C@Pm9�g�cTp�&\+�FE�l��@�����+H�:�Ԟ{�T�DD� �5$��TY��H-a�Ȥ�¢����K��4���Mm&�� ��6vԤXڮ*�"�@}2���oT�o�HAgcǊ���H�
6� 