BZh91AY&SY���( �߀Py���������P��r����r��#DƦ�z$ �h@F����hD���      
=M�2yOP4   d �&M4�dd�т0�F� *JMS٥O�����<L�ښh�@M��]"W	"Y_1�b���%Z��a�SIXHe5��͸rXgK2CGUQ�!H��^�]~��͏6φ�7ӢqM4ҟ�s�#f)ǻ��]6V� ���Ѕm��x׺y��F��-�����@Y�R4�+��@���|B���VID�k�`k���Lq����&����o��6�7W�`x��3��Ү:�o�w,���`jΣq��\��)1�~%�5�fw�A�:�Kieh[Ma0Θ𠨅���5�d�XF��� �D�5+I�I��I1laH�;��FU,�q^���ZlR�AˊIZ�{%.>�c4Ƅ�AVx�\w43#��M�z���{�j�-zAdU8�L����W:����'��ZS'��Kùf8N#xlcc��m�4�w6��z���G*��T�K_%#ÒQa2�H�$o�ܳ&�b�RC)m���A�T�Z�A@�5�K56��L�j���S���k�n^0�	�!���$,�:��(=�[�z!͓9�zB����*L������,)�����[�ՒG��џd��}���8�#�,������^f�|�����R�Z=��X����I>�"�ޑ������/JtP����)��磺�,{Z;d����-|G!���䦍C�b�f��@��b`��7�X�/�2�l�83���t3�a��i�KAVl_Ѵ�õ_@ȭ������Z`���>����%��Zm[:��#���F�u�6��tL�=��1�\�.p)���vY����DCJ��U��eI�!H�s���tTj��A��==�(��aԮʣ;�.&Zح�k�U�l0��쮶�k�`(��PE�;��2BB4�]"�+���`�dF�|�
Y��ݔiy�Ĭ��sH�p��2|�D�H����r2d�,~G=�m��+��Q)���x�V��:F���R�]��1.<�NF.�cA�48`r�����8pZ��_��b�Y�|[��`�|���#'>�����+�*α�"b�]����clD�!�7$9��`p�2iB�9������&c_�o��RR=+|l�JE�[n����Xsw�t�߃��o�F�0p�N���.�p�!{��P