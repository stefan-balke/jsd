BZh91AY&SY�*N 6_�Px���������P>�gq�aƍ4	B���{B���4��a44�@OSA�hFF�L��4� @�!���4����M�"=M �  ��9�14L�2da0M4����$Hi�	��z(�F@ �SjzL���! TH$�?���9	yBZ&�`QB������
�.�&��"��AyC��o���տ��{3�pj�����P/^F';E�,"`����,��S���{�ʗȡ���F|��h4���+9ϸF+S��4 �~9�A�\���T���$�a���
�QAE܆�Nh���f�곂B�mW3�L�[�l�-q� ܃�;^�L��,��e��ObfќY<(�.2�mwVq�#)+;Q��.Ա �BB�i\Q�L�&AZB�Q���;5!���L�ITh��iCj�*�Ր�a�X̴��7e3Y����lcc��m�4(C����
Kw�P��D�D�]����j�7�U��`V#��Ȱ�H�2�Z�h�cE�|��*��T�ωWfv���by1@�HFWM����a�9�k{v��Ʒ<%���xqW�tr��&3�
D�y�M"*���J� ����S��m!������8<�\�+PQ�&�
�k���|�[zKϚ����Y��l*(2`I��f��d|Kv��4	V��ut691k;5�5�B(K�����B`qhPj`k9�1V!<{Hl��83����Y�ěLC�E[B�^�� �~m���4��AS�ǀ~
�֘0]2�b��:*�Ϊ���x �mP�I�c�>��ʬ�B���@�ퟆ�K�:�L[��d���*l�-��%ܐъ��-���q���+�6�e�4�,K�*04ZS��+�L�	�,��Ac^G�;�,HHF���$P,�25�\:P�4CE����M��z�!=���qS����Hb>r�X>�L� ���G�bs��PЙN���$�� �M ����&)�zVb�Y�.�]�P�(6��q�2C��"c���(�Tfܸb*�+xaz��i$�N�
o5�J�|�A�3�`52&(]��	�1u�0����ާͤc�y`ni0=����X^��)�r�i� �|��;k��R����8F
���a�rE8P��*N