BZh91AY&SY�Bӷ D߀Px����������P^�s��tt�M&�6ML��� �CL J�j���4h   �  �������=M��z@ 4� � �`�2��*I��ĞB4���&�2h M15/��PKI$�He"Y
���%\�?�@^�1�������V"#�0$`�b��`&CW�ѵ�mi���[�j͍W���J'�s�tit�����i��.TN���?rƿ�]���ob�(�ME���s(�m��,L���v�8U�t�D�k� x`q0쥹�z-��'6��q�h5�8��6tf#�j��$m\S[�p�#sU-��L�M��Dp�!��ӿ1��Z�ŀ�l��)qiڋe,�I|R�+$�mU��n�hJ,�҆i�́�b���F�k�¬:+"D�}�!�#�vHTH�et[.�!��j�b\�.Y0(�R��9)���Q��{�_sl�V�@�(����0�r��q�����jJ��jh����PI���$
JIRE��&eXp�-$,\1(cq%����	cx��$B"��Ր��2�d�q�C.�E�a��g9��8(}�����M3�X�A?3�[�y#�b�a��\Ub�����������]<;go���]�;�G�A����Oy����&A�Yt.��k/���8r�w0��Ft���a%;�7�vK�"����'uF���"�z��u����r�f�Z-�Ŧ�U0)�8�r�,��Tf�����´��Cc<	ר�ی�@�"��`ټ��ȯḪ��;C9�X�ws�y�|9��(<�K�tue.�z���,�l�	A�@���cDa
��A$����=m�ͪw�,U����q�Y�;:7ƥ�\ٍ�N~��>�Q���W����C�ld[i���溋�fcj���Z�I&����:�8@�͠W�T=B�(���NaVU_|�	uF'��_�e���yz"V���c��M��ҹi/?��z��Mqa��{��fmr��F�D�]o+��t�3*4��[��f^^��42v>g1֞lM0*�i�9r\�S���h�\[W*g�܈�Ͷ�)��M������<�
3r�-g��R���X�sh�q�J;*����ͷ2�Fdö�g��*JOJ�=�抇�NK�tY�u�_US��e�7�L��ՋDձ��rE8P��Bӷ