BZh91AY&SY�T6M ߀Py���������P�p��A�U J$��=L��O
i�4�6��A�h i��
���&L@`� ���"b! ɐ�  4 �&M4�dd�т0�F� *I2)�L��D��'���L�S���Sb�%vBKI�$h�ҢL�����VM�'��΢d��e�T���*���C!�1$����+̆O[������mݻd���I�|�XeID�s�w���2v����j�M{{w�m8V1%��~�ʻ�3��a�����6vi�FP���X����ѱ���(�7V���I%k�ŕę��+�-�0n�m(��^>J���f"���9��¨*�w�L�ØɁtC�I4�]���qQ\e5��`χ]fn9�c�Z^f �fl$�	�:�d�X���(��E�	&��Qf�@��4p�ى��J�&U�;���� Z¯i^M&d�jMA��U�c��R���U2B���z	:�x*�&R`ڮ�)!Jɢ�QR�FU�q5^!&��óJ�e�3zצ����	,j�KF�y�tED]�U``"I;]b����G,Ԕ�{tMM6��0-fD�*eI�T��ťe�嫘�%�D�LĒ$���$�TPP!,uM�@5�ˡ4�s�+�`�Q��)�(J4<�}�TR��
!�.��M��ɢ�����P�5x8h*���!���1�sLc��3��R7Դ�*g{d�(O�vwu�'��}��O���j�T'�Z7���s��`�)��Rr�~���N�L��ӲI��Fi'�O�rӡ��T:'�^QKRc�ptأ�ֈ�B9��(�����ҥ��h�.�v�S�p�l��y�r����v���u<�\�VS��h�5z�"��s0��43گp�WV�����.�0��f[$���&�	�&/�ݷd�J�9�e��M�㿥��6˿g��iM�=�jB���匠�q'T��dI���#���Acd䨇6s�OW��*;��U�Ts��󛶴2�&jW9*%��3�U��{d����d2.��FE�V3�ֲ�Z�~+bFFYӥM{�^-Q���Z�������FO��J���'�ڋ�nyg��)<{u<nW���w��pv���9_m��7�%3�<cFP��󍤨���ǨM��驣��q�كauT�p�gK�2�aV����l����ؙ�3�u�F�^�4_2�*կ�fה��nl�5KC���5q24�D�1��&p�uxK�*F�ߝt�tT��ڳ��q�o&M�q7e)�����S�i��H*�������H�
��ɠ