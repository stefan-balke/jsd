BZh91AY&SY��� 
_�Px����������`�y�s4 �Ԛ4�IF�mhj�M@  �@&�(��	�h  &C��b�LFCC �#	5i55OzJ4�{T�=O��� ���s F	�0M`�L$� &#)��j4�OSM F��W���E��!�I,�{��W=)?ʁ���Kg��p�� ��2��te�UIj�g���}���~׋��ǝ]�6c�fLL�L�������a�q�,�7���9�͞˕b�b����o{�yS�̊�IJ
�.�F����gD}Ȍ�"jp9��,��77�W[������b�u
���r")�p䐣
�>�-�K�����pe�d&�0������i�z��_x�O$EL�9��C(T�T�(M%$���q7����#��+[F�F���9�{{��s[����ȆA6�ST�Q֡��	�`�1m�Dr�h�keR͘� 2�Y����탐0�)�V"�@��\��w��'m��-��UR
�������q.�))޴ْ�U��e��t��r�a�*3Vȷo.���I��0<��\c[�� ��ó�Z�ޞA[��sa^3P�-u�52 
,�I��7�XR@T"U`,�S3#GBr��
�a)A�y4�ݰ���v�ƒ(���w�ko��F�^#mj��^]�VU&*�H�:�h��U�5���+��@��"QGL�p{6O����� �],��*��Ab�tj�ū"�E�)V;�-0֔R"�kk�1,։H:)��I�Rh͖S;gʒ�E�o7��}��"Y)�r��0qXƋ���Uً����Wa���X}�`&=�)x>}C�DJF"��]�j�aB�@����dlI��/�$0L\c��vp��8o$^�a���������������>Q����R�RK���?��M�v��r��4.���!��=��QGy�ߒ;�����`�t;�YT�}-�ۢ�u0E0u$�/���3R�W�B�u�	��sn�(X����<��2s� ׸|�r+�?{����%�Wyޓ��a���Ը�'�ɋ
R�Һ:�/n<��p�*4���'��jХ9q�1���?�ʧ0�V2��]����4�vYc���P�6ah�(OW��l;����7�gv�-�(k^j���cj��_+R�:��"��C��*�d>Ҩ�C@�1��./���.���dD����v�ޘ��wB��^)��Z�|<=Y��c��~qir���r�S���x��HJ񍈨�R�x�'&�^�{�M���bpv�g�b�����r��V�kE��M��͂�z�kLm�9���K�՟G����Yk8�5U,�T���6|�d�yi���!#@�RN
���d���FI�r�Y�(�����Fˢ�\,z�i���T�,�~tڨoQQ4jf��ܑN$.�_�@