BZh91AY&SY�� t_�Px���������P�<�!�� Tښ4�i�	��d�@i�ёDL�  44� 			O&�OS���� �?T� 0�b`LM&L�LM2100Q&����&CM5 F�yMy]ЇҀQ$�AȐ��N��S`�q&��S_#�v���K1��� h�������ݿ���{������c�=B��2�����7n�Y�l��S�m�y�l��|��c����4�J03#3Q��lԣbq���k�m�-J�^�1���v�!�V���B/*�����1e"�i�n��-�jӤ%31)�/ �q��i�����-���M�,aN���Iz_թW�_ �h��������d��hR��r�2ɮa�-� 0ə�p�\�!�YT�£�R饄�I�w-FK
J�H� $%C� JO*���k�eAk�Q��K8�����D&���*$�Z�54��]�Z�t�F61���m������~���r�@;�։R�-b쬌\�^F�#w�:�+d\�X��)xF:��\e���-�#\4K)�3��t�d������K�g�����?x0	��F<.0�m"��Pp�v2��uqaW��о3J��;;SvՖYc�K����(��Ly����������Ȥ6i�mѵ2%H�m�#�l�}#�PŇDw%���Ĺԣ���+�ij%�F���T�)R[����%E��<DN6�]vk\��#��y�o&��dE���:�����ܘ!��X�kX�*ȟ�8alC�>Y��>�1)���nB��:}�Q<��60{["�iT�_C�~+o�HsءB��G�d9��W��I�Q��Z���]eaOn[��)�*Ы��|[�?f�1d��
)��O~�Jv�}ݜ7�a�5��U7_�=ݎ�0�]�O\ɕ�v�^��8��J���Yu&k-u�5,�Z�n�PGd�\��)bBB4r]"�\��2�k,�р�L%��)��a�p�NV�����+_~0��TC¾����r����X�ҷzzMi�K���Ƚd	��L9�I���ʊ��3/t��|�>����M�K��b��id*�i�ǅ8�Kv�zu!vs�-��b�p^[���9�(��r%�.4&)�N?5���,0�#�m���,��I�k��!��w�嘉C�c����#!c�u�k�o�C��	��rŷ���Z`�I0��]�	���)�|�?H