BZh91AY&SY0�� g߀Px����������`<�B ��d ���24�4z� 2  �  `�1 �&	�!��L��`�1 �&	�!��L���B	(�@�j�  i 9�#� �&���0F&$&�&(�#M)�OTy��S�@ �OF����$����- D>�7�:: �A��@ċL������}�F�B�2�!!��Rr�J���zL��}϶��s�jS��3�����'!�sL�y}/���<��M�WӮc������J�x�?kăҐ���/���T�t�T��s�/����.x�NkP�qS6NG.G{�Đ�i@IT-��ir����ta"R�7Ч�����;�*�	&�1ݗ���NW�x\.y��_�dE`/2������A~CgW��c"GT��.ٹ\1�b�)uZꋣ���������|��f�f餸�6e�oriᣍF�KV��lm����Fj����8�7�Zo[�u�Mh�zPO�BN1jEM�1a�2�5�����Z֙��ŋ2R���k�jͲUك�0��4���n��6��B�+�K�.��=[�V�I0��5�%���^渵Ӛ|��w��d��[�#N���T��m���m��IA�f|C����H�B�OߢT�Kb,i��66=D��J(�j�nI��Y	�F29d5PtB2�$xف�T�"�T!��� lm!�^�cL���Ǯ�;�k�����<:%�2�"/!L���eء�����~]������wwwX�mm�H�5)DB�Y�����8B�7��B�kI/`h7s���p|������@b�O�;�nxk����}4����y�jK�"�����G�e�ʡT���ּd���f����v�<KqI<h��^ZcI��]g�� ��<,��=�+��$���Ɨbh+�!�\Lf*ʟ;;��߼����I�Ї(�7j	�z�� �]�����PP��;�����>E ėOM�d��IF�E����D,膋�4,�^�b�``��	���}0������$��r� �/=Ap��0�XX8�����Lė�Q������UA�0*K�
���0��'3 ��3wI�"b��ђ�A�V:$# �I���Yg����v�,ҠM��2H�[��r�-�ԉ�� �G���}�֔@z{dfs�M��{ÔhL���6�I$��)&������IdIL��h*o8�H��X4��i�6�!�D"c�Kh�Pf��p��4ے16�EI�Rz.�($�.�f�H^5�\�m��$��[ۤ��D�A����K��e�{23i4y>�Xhh3IH���q`2D��~���'2�ko�̍ �0hQ���rE8P�0��