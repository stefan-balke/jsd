BZh91AY&SY�K�� �߀Px���������P�q��;����$�4jc!3TM��CLЃ&� � �        �(&���S���6P?T�4 ��`LM&L�LM2100I
e4ђ���S���z4�y � 4=OI���đ[�%�����"�W���*�2=��U�R�=�UU�� �hXL�I����$b 4?F㷆�3���|��_6z#HV���#ǳ��wwEևաC&�F�uUl��Be����p��C��՚.3��:�C�SP��,
�lT�g궈�ɤ�PY�]R����E�PB����c����דİj4��G���=�!E�6�uR5��g4�kj�=����`��ߛU�e��`֬�Ɣ��3s�4b�F)Rk��%�%��$D4�J®,d�Ø1�*���LʉUR�&I��d�G�N.��l�QG�s
,� �U��ep�
�A�P,�c��w�̺8D�����bi&+E�i�Cx���7���hixz�>���.��w&����>�5X�3{��b��tT¢��S*Hi�D�du(^�Pؽ�7K1��(�N�T�J�Tj���=���ܱ�����ӑ�������v����<y+4����t"~�p_�]����cE�3�����nj\�bZ�r�>�]l��<�*! ��=����=Q���R4��
��6N��m�ژ7��5�xO��r���L�8�ԙ�����K9^�����3���J�-N%�gu,��x����M����Z)��j0�l�X�ZcsV@����q@֘��M����v�Z�r2lZY��m��Мm,q�4��F� m�dPY�T�~��/�2�R�y������;:��86�afܢ�E�B�3wt+T	���F�b���h�H猍-�ф8�wf�u�ſD2$��Jkw:/���F�^uv�t.�f�e��5�q�1�!������ jXX���XD�;^(�"b>�(�C7g`�Ռ2b-Q��dE�KX��m�����rڇc�0)�߭%ԏ��y��ng��.7�n�S�9�cӅyͪ�L����5�+�k�GQJ(���!��<�M,ݏC��Y�p�N�3��1�g�Ƒ�#s%6��q&V��M�)�ݝٱ���Ÿut2B��p�cY% �d�È�uDxF# �~*i�O0~���"�}�I�2L���S��C�f�,���g>��UO<���c�5����la�rE8P��K��