BZh91AY&SY˿�� s߀Px���������P~q�1�  ��iOQ�0�@0���Lsbh0�2d��`�i���!�Jd�I4��=�T��� �z���sbh0�2d��`�i���!�*H�M���4(i�h4  �'3����Ld�r%������v�=��U�I0K/S��5U�`�kTL�@�A�Q2pAf�+�iǻ)�ฮ+�erF�����$~����ѕ��Sr������xj����y:|R��=�����.d�
�	�L�i
 ND�'2(=m_0I|QJ��	#T��F�V�\0�CI��,�I��~~��P� ��!k_c�/7c{O�4�{Ւ�D�;���QO�E.rᶑ���%A���F8=⁅ڦ��HBf��H��X�V
�����1��E��R� Ű`�2i8�pdA�7��qy;�6�8�J
d�V��YE-k��ݭ�L'7ڛ����g#��Jz���f�2w�Q!	KrI$�P��^���#��4���dr�n��q
��x��AܐbQf�i��n�#̊��XfA�̒�{� �Pe;�+���8��#}^�u`�����p`,���q�喢3Tk%	��Y?s9OA����D�ь[��@'@�v�^��忾w�g�o����*��-�F��-��)��)heq��0��?�?��ROw��({���On&)N4:��y�B:����C�_����R�����J���t�Υ�)h�6�vT�S�vʒ)����N�q64q��&#�����C PE[F�O�Q�z�a�]z��GK[�b�2_��=��=�'��:����nq��e�v0Y�(���D�]����)��0|������s{Y��M���׶o�X�o$�p9�іYx���GKt訓~|C�����+��ቱ��4f��vچ:�U��5��;$�ab��ȹ���,u��Cغ����_
qS5a�&j������s8�t�=q+�[��w;LE4z��u#��3ף��,;�~K�܏I�4x��9�Q)����3^
�Fm�:�C��I���w5�4��dk�d���)�غ�C*�W�6���nLT��˝2�e����ٰ��^���b6^Ye86ͧ2��ŉ�z�.g�����n��YB�&����T������)����溇vnSc(n�YǕ�疪����s�?*h�oQQ5�xj��rE8P�˿��