BZh91AY&SY���� ._�Px���������P>:"�4hI!6��A�A2i�Ѧ�@� �M�9�14L�2da0M4����%2D�)�4��i�h��  `LM&L�LM2100	�1G�m"b15��� ѧ�H�5�@=�	�@Y$@����A��#�*Ф��2My����x�B�4+&Y�	��ԤC"D���da�y\�3����;���D����X�\+(�y���N�Ց%G��9��Dϝ�s���G�+"��X���_y����&D�M��
�1\oc���q�1�XѦf��]O8)*�|e�Ġt�i��^��˹�x�ق:��ԍ�
�Y���Mq1;��8<3$X|[��g�h!��F�N@��&.�⨩�X��U�T�2A5X����M5
�Z&H����,2AL�c.s��/��������Y�Er�@�_(2�#NL_4�
��U)�i��a�����I$�
c;܇g�<3��i�$�Wߑˑ�[�RЫ)!	Cm!
��''Ib��
� �"DT��e/2X�5��d�eM�3U����|�f�AŠ#>�LƫW4M%�Y�:|)l|����<v_���ILٳg({0�4��l�e�$.�v�V^��v��I����d p6r�P(�80�"Z����_c�IU�4��K*�i�O��F��d)���{�Y%��O
�[]L�n�g���Y�6�B]��&Pɇ�0��W�+
U�s=Uև<�-]�bdS�0�W�~ b�V��.2S	v���)�I�� ̒�G
�����v{ɑ�P�IM7��qE�0S<	���a˸6~�=��X&��d�WURy
�[-�dXX�:���v���+�Sa��2ı-�X�2(��3�-ϊr���-����HPb�N�ccQ�� �\'$u�Xs�"�D4T>��Q6DX�o�}:!=���r���N�R$w�#�{v��$q���#���O�>��)�{bHO��l@����t� �*�LJd7Ǆ�y���(6��3���G����#B�3ݦ�V[�K���bu	�=W�(
�� �20X�����\[^�d���N���
*�Y3�L��cH���bni0=��a���R,m�/*�2D����ב�R�,��B��~f���H�
�� 