BZh91AY&SY��O _�Px���������`_��   j�F�SC��2h!�#M��4�&E$ѣF�Q���@ 4 9�14L�2da0M4����%=%51Sj��h @  4 ���a2dɑ��4�# C � SMOL�LM�<H4h �	�/&�@@	*J�H���~��Ą}aZ�H&��_1�m��4�hVf����9����oᣣF�lp������v�oYk9+����1��	��2�y�8�/���E�����sڕZ12�����7q.��NoL357�w�6Ӓ�̲'�Pc ��c��Db���B[3Ҁ%`̃�KR����m��[���>E� �Lwj���|"����>����sD��2�r�^T�jJ]�g�0�a��@s2(�N7�*J�t�*��+�0�B�,(&L��S9�g�YmŔ�mAA5X@�h��l`bg02�æn\bhm�V^p �P �
�Y{�H�C@�P��x'�[.����� �Gq,�P���%*��]�2Rhf���Ty��h�T�rj�Zʠ`+&���sQ�Tl���
��C
�2�	��vw69��PbD@�cc�(1I[��Be��x�:��.�UhB��v�w�F\,)���.Y&Y��K�#�s��ܲq$1��"�Ȥ�j\Ga"f�����; W]0&W[��Y�a`�k�o;�5@�Z�m.��8KMS��6��:���Sx�"��@��>�7��5�Z����Dtu����޲"
�6�zM�����$L�A��m�����=�܅��i� ���o�q��)����������2�^}�U�H4b�GցA3[R��Y	��%���<�u��	V�͡i����:r/,�Y�.�kT�!mb7&�3�D���JH�3����ϟ�
��(ć�7iz���z���T�B]�x|?�c�`��A���G-QѾ��ͧa2U��Y�S�լ���ɜ����n�/��NU05$��-M
*���ʵ�f�hh�h`Mv$�a�G9^��6h����Oj�	�
s2
�s�rQ���^@9�P"A2J�Ȃ ���"��Uf���H��*��&Ȁ����b�N4���F����ْg����=�LB ���i�K�C�1�2�Q�,H>p0���o"@b3�qc�u��x�t�8��i�9yI"C�g~��Xf�M�
���s���i'P���?)D���C��g�qB�C����$��t��T@�$H�X)v4��^���ĺ�7�4��@�XԳ�B�H�f����_#b��,��BC������H�
�0��