BZh91AY&SY��ܦ S_�Px���������`?-�eh�;� �<%
j��覙?Q44��L�M�L�� ښ=M �@� ��5'���� @ 4h  ����L��     sbh0�2d��`�i���!�*H� M2'�=4)�H����bM<MO)��B�`-$���3�B����WlH|m�%Ԇ ��|�U{�IJ��P��yRI�@G��f�=�Q�x���ӳ��7i��MN�K�g1�慵N����{&�ڲ�[bR.FE@��Y�V7vU\5�)����D��9�^Vl�fm
¶�ֻL����way��Wy#d�Z�A���/��347�7���E�z�o���������s���J����>�C	��;B<n��ӱ)�̕$2[i�&��N����u
��l�	�K��sU/�e�VV٦�
��Q�M��mK&�E����RTFPEk:B��S�83U�^�ccXCT�`���At��/WwK(���fJă���l���r�db�RC�����sͦie/h.-U�U�*Ca��ы�4��+2�k�0E9���(��M��N�� �Ӷm\���ՙ*&	��e%*���[v,�Łg�B � "I�����[��M1�S���N\��P��Ia)��F�6�T��h-N"@T�:�D�aF���{��qfn�r�T�k�r�T�+߱i���A�P�5؝y�����)��M{F�jrӈvi� }C�(�9�(�s��a�Vk�04`��s8�B���?7зĹL���t��<����D���б���p-�q��0=e-<�'�����G?<�Ϥ��d����8S�㑊S��%��g�jqb}�ΖY�g�$��ľYg��Q���:��}J�R��h�F�v��E1��T�5AgЌ
��w�;K�ؿ���튲�M�W�JH�pb�����^Ѹ�zg#�C|�,b���?����u�+�OR���ǇvQ����b��qQ���ʹ>�}���[��{zr6|Z8���M[g]ŋl�.�Z�e�^=��l�Q#�]��x��Q�w����Uy����#%��L0uZ�^ۘI#Z����Rȹ���+`����O�ldc����SxR��$�P�� 
3k{x���+�=@�:6�{B�G���ϻk�aa��Y���S�)7<����U�w��k���*(�,��<��y��n���K��4���3i��V�N��P��׌mr6s����yv��&w����]�ݛC�f�WF ɮ�U����֩hv19�ѧB�y�G��ү2�M���|jF�s��RTO:��;���\��u�L���ggm�n���vLs��S&���EDӰnA�rE8P���ܦ