BZh91AY&SY�{� J_�Px���������PXo;�C:�4��Q&�52����@mM�@F�!�A*�M
���     		��D��d�  ��A�ɓ&F�L�LD�&�=F��T���M&��j ��F��վ�>�IXB�( {����H��hT1+	2����f�7X�4,�d�	���Q #)C��8w���[#6�q>��v1�3ƚe���]mf�-�I����C|��x���ܢc|"`���È8�(�%�+rbِGs�"Ү�iwϼF���zf$
���@�k4�$��������J!&�1���A�� ��>-j2��(*���M��m����&� p�mwF�ƨ�]�釉��'�M.G�zQ�1�+XAb����Ș͐�l'�%6ǖ��i���[�L�e�UK+X֖=���"%�Fv��,/f�jJ�B�RR�Vb����s���,Uˈ�����5�Q���o[m���P�o����%��#�
I�w(�(��l�TE�т5cu����Y#M��KD�.FXda�腴QA@�5Ƶt ���bӹ���i���qMw��̠Р�4���՘`�Njj�;�_��3�9ZG�s�HԆ����X��5�T��0�Z����YA2_�t��޻���=���K��XHq�h�^#C (�	�Rl��I�)D��*���E���@�����|��Bd3#a���Yn3줞�±��l�M�E%�;��Pnd"��a�D�Cc�Іu�5�R��R<Y�](p3�ȸԴs�6�	Ŋ9�_�~ k�F��^YLP%����H�dIy�#�Q�vW���L�*����K��F�_	�0ҰRM�:��Y��)*=@���+� �v�kφ�4b�4�����gxE{G��e@����b�y�p��0���� �n������@ Q��A �bBB0=��0����3�31��"*@"l`�؏��ݷ!/1ԉ��G�P)G�U=l>�F��;< ���z��g���F������I�a4>���>}�V	�ġ�`^v�ƀ�\�1
��q�!�p�0A��fTf[��U�W �j3�E��Rz0�PJ�P@̌V!�jp(лE�놗"���"�JE���i��o���&�ă���0``�����ZH��8�z[_�Щt��̰�d0hZ19�1w$S�	�
0