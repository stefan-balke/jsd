BZh91AY&SY���� _�Py���������Pr @�h	DS�S�Sz��=P�Q�@  ��2b10d�2 h�00	L��MM5 =O
z���  h 2dɈ��	�����$H�FI�O4�I�==P h4�4�S14�ސ�BE��?�r3��hR
b&�b�fۃ�`+��`e�5�-��L^�&�|{5�ֶ"� ���>n�ʡ�K�b���ҵ�
���Q9���-��y3O��q���~RE���A'I҆��a��#���	"��'4�r���[W)h�
�O�@���c���s��E� �><,�Kq��T�DJۨ�	DG���a�3�~�a��QRv՗b���JXj����խ�+��/JWC�flWM��Lk�7T�`$^�0��2���(hE�qE��%̣#,�d�QQ_,�$&������%ĒI(@�o�퇂b969d�������e~-@��'	(�	
F�ͤL̤�)5nCIa����HH j6�<Xcas^9����#�%{���/W�������q1�+,k�g����I�L�B�_=���(�U��4\�JQV�l�D9��q&'�C�WsG�!��}��B�
�$H��̎>E�2�R^~ʥ�#�:5�J�Dͬk�aLi5�P=�l�ْO=U��Q`�4q��Р��E	s卭Q��1ni(>���+
UQ��Jއ>|���b CC�J-�B�^����=w{N0�.4*C��P�ӄ<��)"��ahLjmCQ�l�a�^�d.�!����٫qE�0S89A�}3�CT�Q��!��bID`0��V,^�ݡ4-!,ZH�v��v ��W�>��M)��X��Q��0��9����h� ��W:�*��llh�X�T1	�5���2��Ҡ�l��^;Ov�'��Dt��0>�Hb=%�}��a� ^�5�Wf�4P?Pj+�t��Ē2��h�0f~��,D��UŎ��dad�P�Nh�q"��D��J�Ͳ7�^�XEo�q7ZE��X(��߼���P@Ő�̘^56�V�! ������J�b�)���=�6�K�79�.`jD��R��H�f��6���5��'�������@����"�(HDV���