BZh91AY&SY\&wX �߀Px����������P�wZi;��Pt�=MI��ơ��2h@���di��OP�@ ���)�	=E=&4�L����D  �9�#� �&���0F&$ ��&M��L��4h ��R�`��PE�X�����c�zK�*hRM%4��5���n)��B�E�8*������e�|��i����W�wY��Y���G�+P�Ө�so|�6�Ք�ݠ,Yh�	)xz$��KY����4�%���[�X�.Zd:a�Azl6))��^3�A���zf�"2ƜV�A�����/҆��2Q*����6����8� P�>=K�6 �S�4f#T�s�* ]�f߂����U�Nhi�]���Y~�M1��(��nUb�Tu����5�:a!b캈�.�K$��B���U��ݰ�,j�0֑ū�
h���Ņ0M]��PX�Q._8dv!�T[+}ܚ@DV��DU���Ŭ����4����:KTA|Df۝�o����+]lګ��T�)��&�P,̸��!	KJI$�@C�CWv䍜�NY *�i�����&TB�u��&�D��CLbQFҒfR�H��i�q((���02����@�o�}�	PDc�g����ѕ�_N96��@���2��Rr�{fP8�z*`VX�B�\?[����U��N��6Ng6���뀊��*����o��q��>܂α���!!q���;�

�d�@���	�ҾC3ڒ�����$}�3>T
$͌K�Z��y��c �ȳ�I�@�UYm46�� �u�.+j��\��� e�&撂[�0k�q6��3�� LGV�#Lc�2�\�ϘVq� �m���B]��w��y(�::(f�Mz�#}h��W�3�H�:!��M7۞``��I���OL3�ezr�Ԓ6�z��@8μ����N�vkC@ ӱ${��7��?S���@`VFԨ00&���U���	! @Hߒ��z
FƠ=��AP�dobT�H�D
M�Zd@EE�2Gv�'��RGr&10B��BG�����b\hX"@o���a�����1�Ƅʺa��r�)4;���"��<�V��Q`t�����Ci�7n!�.�D"c�<���N�Sf���M̡�6]˖��:�z�"!&d2f����/�O�Im,�_i �����S�D�h^�*�.Ƒ��ӑ���{�6����$Vk\�H1� ۜ�mͯ#�R������B�
��w$S�	�gu�