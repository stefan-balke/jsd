BZh91AY&SY>]� Q߀Px���������P>]��.8�SJ J$�O� zS�yF�0�i� i��h!�i  h     *x�"&�j	�h#0FC 	� � �`�2��H�$����6�Se4�4 4'��LH{�
@`J���(��P��4!����~�����\2�!41�@�1�L`F�n�Z���0Sed���B��'�# �>=�����!P����ǋ���J��pt�ݘrc~3,2ƣ`�1���/����(J��>1[s
ڰ��D�6�]�csj�md!b �����>V!I� �LG�.�U2�	Tw��(Ѽ4ϪV����wԞ2�"0h�d�eA'��d�α (�AD`Uh�;�)}ny�т���DV��;�VZ��
�TZ�MC:��%��T�-�W��f�^,��U�D#Z�(�
R��Ѐ�E�� �*�,��\Z�U�Hr�!�Y�61����m�1p�:;C�Iw�8�
ǹ�l��BF�!J���i�T���K�@�m�%A"�4\"F`�� @@�5̵z��%I5�hzY��e�jLWF�3�&!O^���=�	d��n^s������\�[���9Hh�"�ҥs�l�&�h�@SS���f�ƃ� �A�`o}�,8�@�Brܾx�B����/:z�hə�*�V�M�a�@������O]U��Z�Si��l-
&B(K��Ѫ(09�3�D��☖���ŝ�yu2Z�B4'Jsf
���W m.6)�}I����i�j`��d��H�::��g����О�/m��:4�4���z�	��^�8��'G�  #�`=��xiʆ�k&$��܀��z�h�-�>��:�"ķFD�[EjcZUͬx��lɎ������A�(�@���\:L,M�`�J�"l��M���'�g�]Ȁ�w%�"�z�C�~n���@>���7r�l;�>�4&Sy�u�����ߢ �L��\X�o.�]�P�(6��3���c
8D��HШ�,��U�V���Y��X�BjOU�� *;�@�#�`59J5-��Ak=%%�l�r�.�/SH���r9L[����L503	3W�EM�D�7@[�6�抖��fF�q�������"�(H.� 