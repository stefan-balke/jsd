BZh91AY&SY{��p /߀Px����������`?؀� j��5=	��M6� @h 4  *�y@�T�z�2@�b@0`�1 �&	�!��L���B�A���4�   9�#� �&���0F&$41L='�=OЧ����52��܀I!Q$+���ϤO8ؿf%9 ��HbT  �M|�}p/�"�X2�G&��D,�����]��o�6K��L
 �� ��!N�R!I>+����x�]\E���S�[�e��9h��b�Y�$|G��>wV��ai��2� Ȟ*/5�
M-Y��rA�b�:���4!T1-K�����B	M�_L���#��t 0c��н��Aܧ��E�<�����g�&p+�+�ʤ��2����b7�t�+w>ڔ�oո��N��1(���t,J�GD>�1F�"�5Иʎ�I1�	��u�V�8h���-�����B���d�|�*6��O)��koX�޲�օ���n�<��*�\��8����3�,�|&'��+iLo\X�&����wB��=+u̗VL��&q��&�&j�����ws�xs����3&�4�氐֍'E�]��8'��;�$!/I$�P �y(��öH��cNY1
ߒG.F�8a$`nfJ&f%C�?���u#P����H2�hh�PJ���!�a�h�u� �0���� cI&�w�q�/��J�d�Zx[��}����CĥsM��Նǆ͓0	 �t���D�w��q�%n��<���"]�&(�7�}��/h}c��[�0�Axe=��i͠T`�\�X@��ygJu�_1��$�r`�P�E��|����L!��C��� �-�I<�	V��u-����c)kPhd"(q�-�Q&PKjb[�	o�����J�ļ�fd8��Z^�� ����m� �)C~��+�? /�&�Ĵ�LPU'y�z���^i�( p�A�FI��I�G5�[�v�ꆌӢ��Vҋ`^��/YC���~���,ӎsR �*���p��i��k\�5!��g�!#����; h�N��9@h��;�yiR����g`Nf!XnxM�$�E� �N�6�W�������՛�ju()4T;�&�f�؄�d1� :>�z**g�H��I�����blX" ���g�ay��c�Bex��8XI > ^�E���`4�}�Y��-�[�(6���p�a3�%�Lm�I%�l��F`i׻0��Y�7eF'fd�X
�]N9�0 d\ȉ:�N��Q�[�5-�a �����%~y@�C�1���iy5�[I��A���24��a�\T�6���emx�,��s0�r��.�p� ����