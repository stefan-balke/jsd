BZh91AY&SYd&%N e_�Px����������P~:(!� ���S�=#   �   dɓ��&	�F�!�Jz���G��j4z��4��   2d�b`ɂd ф``$	��&!O$f����j4��Ԟ��&�!� �$�RArB�����f���Z���$��=�m���$��Y�!���9(�"�{��u���?v��v2�WbN��Ԥ�~ھ7n�#'N@\)�U�h1����#����eFX���X����I�7����	�Pf�O)�!Z����&T��ғ���<}V]�0c�w���*mnF�7畚S*��3y���	�����%5�J�ʊ�b��X5s�쿛$�K� ���baVY���cB�S)!5k�'��*X�b�p˘Eeu��B�!D���^�ĬT����o��
a2�E�%����\�<INU�Rґ;���*꧟�&�P^cr5t�(�0�-Ŵ�EsUV �M�7��Dm�%��E�vab�6.SX7��[��ض2�v���2)$�(�3q��J^	-�E�[q9�(�M C��r/�Q|%�*��� Bv]���@���0U�{%�����h��$�C�}~�f�!��d��;Z<��m7 >��ut���(����C �� ���}�x�t��* d �<�@����3^))��>����Q&p`n^VB�!���C��d|��OeU���D;�O6��A����ۄ�5@@8�&���0k�hS��Ja5��y�4'��i��c
��3�^6j
��@}7���E1@P�y������@0����_Q$uYݵ��D-h��e4-_~�
.����9�0��c�[n��.�mh �_-���U�sߪ�Y��F�_����N��.P��a�b:R��̘d�Nf�Xn{&�$�X(G=�L��6&I`=�x��Zɨ�E���T���P�, ����:z��Bz���sD�f�4(?�>~>����8,� u����w�3�����Be~���$�}�lI� c��x�0&|�W�<��\��]�Pm<3�!��x8�!`l�EkÖb�"��,��i'P���e *a" p��FA��
Mq(���Ă���Y�"�K@di�R�i4���LG�AǴ�0h7�"���TIq��qŵ�t�Z�{���n4,�w�rE8P�d&%N