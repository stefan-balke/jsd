BZh91AY&SY���� `_�Px����������`����sx�'� 4hST�򧀦�G��P�  Lh
J hh   h M4E� 2  hh   %=(�
&�� �     0`��`ѐ��&��D�<��d�OM5?SA�Sjh h�hjeSB@��B��%D�E�@��x���Đ����
I�Sk��m��&$"���&�I� Z /}���=�OS�w��ٴd�ZH��*�-k���m�m���l�9����q��CK `�m�'}7�V�]Pd��*���-v_v7G*���05�M�}eV���I���<G�y����"�,H�7����,�$�����3T����wy�v�L�x�%b�R 
 ��b��� "2�h��>Щ�n+�`I2ڹՁm;D*�xW(���]4�U�
BA;�
4�X�"
	dਁ%ܤy�=��-D�j�� ��o`¥��]�,A�4B��
`mV�(����<Z/.&�)���J��K�V�@+]�+�&��*��������ļ��2h&[X��EA���d����x�z1U}�_,��wM�2R$�wVf=���yTƀS��nčF��B:�-�����xf!]���!��HE2Un��������T*��k,!%p���˄��������饁
�1M%=Ĥ
`��a�%�$Ә���R�(FN������.��4���b�)eKi{��$1D�`WE)��%P%	3'O�B� .��Xx���ę.B�M\�GbU!�e��2P���0N7_l�!	Ĩ����;� ���Y&��Q��0�L����2�G�2ۇ�I������b���x�M�t��h�(���� 뙫�n��8�JjD�X��N&P�f��DT��QX��"e%(�!2�X�B1��DĩI|�f��ɺYTZ��i�		D��94�K&52P�%� �0��r�;@i m��)n�����'V����;����֚�s�$#+��1SXr�� |�})W�{���]d���#nῗ-���6!��9��I&�l\:X'M6�iz�)vr� �s��{~!��{�p>A 4S��N�<\b�kB�^yR
i�^C4�$�����  ��34�T
$�l+��4�2�}����A�]�$�J���ʭ��i�Ѡ�Y�8��vImj�( mh[S����.rv(O��iq!�ϝŌ���BcHm	8�P��z�C�A�Hg/3)�ARy���'�@0o�BA �Hd�I$n�>�z��V㼡 �]��Y�[᫐�������̞xi�B�9��@A�&K@8ξڃ�z+Z�٭X,iB8��Q���zG�r��d9��z��
�J9�����M�I$#) @H�ΠD�d��ؐ�Q�&UFA�[	�3���_&�����6D,���.��hI�%0����y�;,�W�`���ꑬ��]��Bg_1�7� @����� ��� 0Pf�'�-@�� ��P� ��t@�]Ĉu�����<����[7b*�+�7dIf7ZE��&����P2H�3)�ge�I��uH.����A�n��	)U#�^#!��ى��Ў���{A� �cLِ�#"�`;�\��5�Z�|���B#����]��BCKC��