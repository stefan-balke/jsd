BZh91AY&SY�e�C �߀Px���������`��U� 2 �M#OH��     �� ��    � ��T�S@      	OI&��L@ �    9�14L�2da0M4����$H"e<CSMOM4�I�#M 4i�jyK�h$��!@T -(>��r0�hRM&���M�|�B�4+cI���9 +"C�����~:�zKSӾ�Zb&f.f{�����.�v}�ޙHP��x�"y�N��!� X��#A��M�	Eb�v�ZÊ9K�ٚ|�x}��E`��d:R/�����^dF%2��M<��o`�V����Y�i9��P�kЏ@k��M�S��V�}%�y@�@��1ٟ˜=��F�v�7����Q��ky%p]-}�k�J���l�}��zV����Z�&��o
�[�CZ!
&x� [�]"nVe1��Sga����)1 ���r)B��E�����݆� �aӦ��'k�s�d��5i[��m!Y�S���$NH|�W��`�	VX�BK$��}���B�f�k�c3��pb���J�PA��l���0P���)��(�j�Z\"�Y�t����yJƈ��rR+9AAQ*^\8eqX�Rc*d5:〹�b��׽�!��������%�o�\�oH[3�ݽN�(�"磌BQD!�� �]WP��]P�;�K�I�H�(�!�^ࣂ����Ȣ6*��%�q��.]��s#��U�s�"b�muP�n�,���[�ě6�k�/�~_��_qm��ը��`���:L�0aRu�s@ɱa�����6��Dvܔ2A���0V�332�Q�8f�]p�@�|Cv������>A�nC@��!!y�����
a�B$���H��}�YȒ��ED��䌙��@������؅4C5�õ�A�YҒxP%Z�n56ݰ����/,jl�P��kTHe�ַ&�3�D������UK�f�އ>���(�'[�5��gH� beن��%1@p*O����M:S���]�����-�i2uCE%4,�^��`�|	���y���^%�����7]�͂����,���k�ɱ,X��ב;��X�����k�\p��KI�H�`P�`�2s4�a�e9F$�U�Pt��
,0A�3��B����P��yN`��0Y��4`�w�TQ0���.�D'���#��7%@���G��s�>�B ������F\�����p=Fఐ�=�`!��su�FA4��Y-���-a[�qӚz=$1�G���dm*3_�!V]��6�"�u	�=z
 EK�8A��\Ax� �P6�[��Ae�H�),!Q�o)s��4�|��N6�Itsp5��i,3W���H���;�^"���ّ�B�
����ܑN$.vP�