BZh91AY&SYr�ܦ �_�Px���������P�s���2j�0�DȚi�����h�m4�� @�U?S�HzA��     ���
���OS�OSj� ?T��� ���a2dɑ��4�# C T�#4�h�&�z2��h�Fjz'��_$W�BZ ��Id+�����O���D�Az��qﾪ�v�J�a�Bh���Q����N�~�#oΌ�y���ͱ�k���O_w��9�f�r�*֡�m��H7�+0_���[� ��ˈ���E�L5h�\��lh�3a+LWpף,��rV��xI�U���LNC9_��^��|i����N�΅&{v�}��#5�18���q��,YXf!T�z��1u~���Wb��Y��3t�&%wL=Gp{&��G��K����d���R��֞
��1�g4�g�lp�!PҬ��H�y*`�DV�*$�R��f8vq-&�%���
3�P�r��T�Y�QB:.,\��/q�k����Tz=!fI�g��u9�lc{6�m �=�l����R]|�B�;ς�R�*�2�k��e$��c��6������R�G��j��
ʊ
�����!T.���Z�����~bH��L�����I��ֲ�g0�,/�E!��Q!e�r�	�	����rF����*��j5�j�l�'���h�@�mՉ1i�jdgȤ?�б��y�[�rqr%�)KC��xqC�|T˞I�֘����S����)�C�w]2�KS{s����)e��XI+nc��0��h<����e82"�xi8�t���w��3�"��4��*�>VsƨpgwK&ɫ�KETR*�5�to32��2+�V�s6��������{}�n�(�<��N�P�zۯ�	!Y�APsbA ��P�/$Fe�M~:8&{�lr�ѯd�X�n7ڮ��ai�7㲴	҅DD��	�2 �n���߁���7h�u��͔��n1�;v[B��.�,@ Q�z�(,A�Ą�b>�Qt��ak3�І���E�2�$Z�ZŲ��2}\�+~<�{gB`)�ѵ%�G��ߙ����Xy}6s8&�_�]G"�S���y�HW�6����q�pCB�h�ߺkf�yڏ*\����b��|(�Ȩ1�+������`g�݅��ht���YS�NE�4����-�Q����`8��L�ۆ��z޻�Ht�w�0�xV�*J��Y��r��p�̜&�(�tY��ۿ��w9�g��ECz��\��G��"�(H9snS 