BZh91AY&SYZf2O �_�Px���������P�wX�d8���T�������h�@6�L#!�@ jy@iOT 4z�  �   Jd�
O�5 �  � � �`�2��H�D�jm�4�=&�~�� �ɢyKɡ'�P�D�,H?��9$�� �B�i)��A&����n�bA�pE�@�Pv�L�M����3_&�^M|�W�RLj&d�M�x�^C����\��5`
F�9BJ^�<l�j�~�g7x�A��3Jai�9�� �5�2�X�1�:v��d�t�BJ�h�
�����5D���|�6�R
���zt�L����>�F���������*ʬ�H�'bj�b����؇X�����-jZҚWW�Rh��#$�e� �� .�q�&L;I|嶨`lE�5�8�+������Ld��ĥ\R��wH�T��ȥF7�h\�v��
C5aY
̹F�D��	���e��wM��9��U$�!'<1��`E�U�R�V�^��Bs�VE::���#�/�A�	�)$�
��\��zb7r�9d����9r7K�Đ�HBQ.e�lHE��RR�YD�����r��h#��"��)������Ƥ!D@�h�{�R�����6�ֹ�
� ��g�ym��AI
]	,o��h��>��Pt������k���h�`�a��_��!m�Ou@L�5T�0g���7�`	�H^{��~�L=��A���^�����n䗟j0�1�>��9���(&b�ּ�bf����� �,�I<h�l��6�g�����5�B]G+T��r�8��WE+
U#�=U�yt��BM� �"�6a`W�|@�n�b�-2_#����!�tթ0`."�6.�H�:�k�vr� Ψh������qE�1S;ɜ�˽1�HBIP�'�x	����DD�x8d�Eݨh�ihA�w ����4z����΁q�i,%�*�$��s9���I4�h0Iǲ�*��llj�!� EC vGDD��b�5��X��E�rG�rΚ�]G*&1>�RR�Iq�;�6�HW��q�F���!�cBex��,$�>p4�����vmdg�KAa�=���V��0
�4��!�p�.������o�U�V��r17�"�u	�	F��J��]""F �j��-����̐���ii��&/ �I�>H�Ƒw�ۤ��b;�8t�CX,5����H�v����&�K-�Y��f0hZ0;m��.�p� ��d�