BZh91AY&SY���� 7_�Px���������P>r*(����JI"��2z��'���SCC@h  h9�14L�2da0M4����%2M)�&ڣ@f�!�z�  � ���a2dɑ��4�# C � @!0@&��Sh� �̚�1&�>)$B��@�@�_��d��*Ф0Sd��?ɶ�_	�W�
�,��D� 56��Nƛ�}���o���{Vz�p�Q#��|�8��8@���#^Z�i�G��l��p��m�*2��c�c�0O3)A��e!�0���f���3
�wNhP�?��1��k+��埼�u	4������E�;�����k���e��E�R)%3�E��XS�S0�3����P�!��P䝓�K��Z�d�����+�rd��6��-		��Yd�QP���8�
`�tw13��$Y�N,�U6rI{��14Q[ݙ�՛�1��N�$�,l�WT��q���m��
"�nC�����rɁS�H���j�ML��U�ClE�	��Rm� V���D�h1�2��! ���3\�`L��/�Q#6�wrN�"y�v؄�N@���I��~]NR$�R�Պ9ʃ���r���R�:����2����i�31#�]�fqA��xԣ�]!�V���A���S�K��� �ݜw	")B�a� ���`ƾ�7��$�Z�H�Ј�qQ�P����e�%d&C6�(��A��rI�@�kk����e�A��E	u��Q�+K�4��&a�)T����7f�<���K��C���B�^�� �������(�cp{~u�\ DG�������[��v�$�6��з���o�U�4S=��pf?-7Y�cVG ����P�k�H�M3���̐��ĳZd��~�ۍ�%�3*GP`fL2b�͆�����o���$����*��#cB�OĔʤT1	͜"�,ADI��y`�<���z��g�K��T�V�$0��3LԐ+/!�keqQ��P,�(�A�d&W��9�ĒO�р1�Gn�-A4L��+���8�Hu�
��[�d�4��i(ًX<b¬.���>�Yu_,�B��Rw��PJ�L��d�F���B��H-a��Sq=$UjDk�R�i�O��{I�� Ӭ��!�L�ڱ,-$�Ì���ב�R�~���B���g}���ܑN$+lc� 