BZh91AY&SY�H�� �߀Px���������`�xu��;pꀠ*�d��z@h ѐ4�L�O@
���@hF��   `LM&L�LM2100		M2Ħ�Q��iF�h=OP  � `LM&L�LM2100I&�LM&��zL&M  zMKȊ�$�cL�K!_����h6!�A�B�1! �
k�͛p<r-�t2� �G���H��>^s�ѿ��<�Z|�ќ�wg'����&�m��'�O�`��f�|�$p��eC���F��f��*]	G4I
�߹Q��������\��;Zm��[�7����9�	�y�V�ӟ�&���fם��I3�?h�E틙D�x&�ᬒF�qC�ӿ��;`�4��m�g`w�Dh��2�n>kg�̥E:��^5��%�r��.(h�KdATE�Җ�̻�9Uf�Y��l����+el�G{,2�3T�����(rega����0DV�r����U�WKhSN�LĈ�	M�A]KD�K.�GA�L��ª�Ba]i1.I��.�\�m�c����2�l03a�1��KAD�:��CU:�#F�Ҡ�v7�(6Ej	bV-@]h2��	��
�[͹�Y�k
3n�6׃-���²Q3U�b�P���FS�.�����lc{�m���C��=�ꤻ���B�i�T�L�b2UP��؛����2.2^d��cj�n��l`輀��i��fUJ�X���a�l�1!� �6~S���~�ߌ��_~��.c�
�6s�IMBbd��]t�jV���:*x��ڢ8�x���7�
��fv vt���JRJ��hU4𺤇�x�N^y禧�����4d���Z6��l�z۵nK����D�L���|u�e�ꙹI<5$��HxF�p|11Jq���L�)jo\�}?!���`��ƛ��0m<4��;6�3T�}-���nU1��(r��J$�X����w���g��u�7-{RP��*��[��o*��1\tp6��K���_����͝r�)!l7�x���]3G�ۛ�h��u�EF8^'
��Ō��)wл�SO�__BY��g߷��!ן\�DX�nh��jVܲ˿��Tk��֐��JC��|£��r��F�M.�i�c�о/���6�6Q�y��W�~e���"\����|�0.A�=�X�HF��fi��Y3�u^엋Tdz���k��'��%tc�!�t:�b)��󉂑��ۘ�s����=�������7*'�v;�#;	!�n��B������6����t���;�����#��U*�WR�)K���E�m0j�&Jp�ѩ2�e��&�,�3/�y�h���!�N�79�1�R����3�Р��r-[��0��Yv������t4�G�ggkq�����Dl�`��c��6���k��g����n-���"�(H�Z܀