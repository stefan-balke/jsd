BZh91AY&SY!��$ ߀Px����������P���@�8�	 ��S�*{Tzei ��� 4M ��M%#@� b �@  H�B��#Q�OP�4�h 4 z&�� �`�2��H�h�F��ѪlhF�6� ��CL��R@>�P�
�B� @�s�v�Ў�Av�#�%��} l�H�hU��!��Rr"Do��[���}����|UUfUW*��QH��w ṵ<�e�[;4 Q��,m��s�:4�{�}��2�#6�� �Ήe���hy@�
�|�� ĤF�s*�2�s��Aj��x�$Uwf��
��V/�� �H�
ҟ�_�H��j\D�L�������9���!j�W2��Q��la
S��IuA���$����\b�kr�Z�Ye�M�=�s��1N2�3!�I��e� �4�%a�� �-�9�H�齢%C�Q%�CI
�+�����B�@/(������D!�)@so.�c)\���8�֭3!C!h!���(yZw�D3�+��+4U��
�g%7;�#JFEV�������Ege��a�܃k��0�"�m���PA�GW�:�.^2L��rIDR�����˚��U�cPư�	.��w!CCp�a)�H�0�Ȃ��BA�5���1$�3{#9D��n(O�B�.�F@�˄���U�����Ֆ�}��@�
oRi@���l�2NOyxn�綸�#6�D����)�Y�$��:2�Z<C�!�n��/�B�9���tj�`2#Q���*'�/��{�T�"�#�$�ȹ��Y��f�R��"�5�n� �a�I�M�V҇sKQ��ͼZ���DX��xZ�L�K�4 �u�`��Z��z�ؾhp3����W��m���N/&sj
����@�����@L�a���� ė$c!��đ�H����$A�3](�B-��-������s�^�g f+�����^��l�S�>���,��M����B�p��26�/Wa�E�����aY���)�JC����i��)	���T��lhrD��"�������\���Hz
����ݵ	�Y��%���4��zO/DT�LV�@�A���E����F��y��xTI$�0$�`1�1׬I^%��>�+��V�0�hLm;3,�Hc
l�a��IpFkە��M����ʩR):��&$�,��A�3�@��D�
L
��P�.-�W]"�$`F�GcH�����h<7q1
��H�֬)�"��{��mf�:���e�"b0hY�L��ܑN$a�	 