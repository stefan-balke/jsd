BZh91AY&SYź� �_�Px���������P���88*���#E6�є�F���d�z�  MA�R        H�����O(�z��SC z� 4���	���dɓ#	�i�F& �"@�6I�"baF��� 4��f.IR@� FJ��w�p�%��hRLbI� =�m�� �hVL��	���
eP�}Pb�w���pV�{���=�&e�A��FB�;_K-�oޱ}lP[L��Zt�7�&�2�>6������	�b�1Ϟ6slO5���L�i)��ᖏI��nx�� J�sB�俠{�(�;��~�t����L���p�����+��:(IdN���N�Si;��-�,��^Qp�Pa��3i��ք顾�T�#4�1�nb31(iU&*��B�z:5lD0�B�x4p�;Jv�Yԣ�J�K0��� 2b�&�����C���P��K:�V��eTW��׽p8�%�/p���T��Y�r�MCc�v�m��Q��v<A�m�)Ԣ v�*T*�/��#)1�u�i\6V�J���(�JqB2@\,�e҃*.� 0�����ěM���Y�m�xq�M��%� TxR��[����3I/T��'>g�4�@�\��q2��k���&Q��K+����Ҍc+�9��z�rA���o����wHe=���
B�u��QP��Ð]x���쯱��{Z2��V�4"�4�	D���aM4��hT=��A�wzI�@�ku���;��fGf���E	ua�D��b�@΁��VI;�3�m�p3���*�����m�43(r�
����߼4.3S	w�����,�U  A��@�H��F���ن`�R��Q�fC"�
-��&��f�l&rs|����]�n'N�D�Z"T!{0��uR�%\,q�2 ��W�}���P}�E�q�"a�9�a��9FD�1 @H��EI�	���D�~D.��vf�.�T�!����D��]��	��i�)��L��R#�I�X9i"]C�ŝ��dL+�/�g
�7���Gq0�$��F �<9���r(�,�A�^
�6�Ӫr�d�4Y�䉏by�A��k�������,N�5'~�*a%�z�V!�jjT8л��4�%�6�)� a)��_;H�����&�� ��n��$Xް*#)"x�x�י��<ʷL���$)���c�����w$S�	[���