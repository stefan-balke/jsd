BZh91AY&SY�] &_�Px���������P>������:Q*~�j4��je=OQ��4=C# A(LE=M����  @  $$D�&��MG������ 4i�`LM&L�LM2100I$�FM4�G��cQ� �#A�'�� ��"��2E����W3��d4*�`L��?H8�tXB�hX�1a�6��� �@�)�t����7l�;=l�z��l������^IJ�l#���
,B�1���?r���U���Ur��,f+��`1dW3˲bL�]�xhiX�f����M�� %C2�g8�2<���-�.����=��f����o	ʹ�5��Ĥ5 t>��F�����	[T#y��,���h�ad<[�AlULEJ!R�E����Syg ���6
D!h��&�aY�0B)�-�W4�gR�F��	j%��ckA�*S;���,Y�бw�� ���7��m�4(C��8|�Im�ʅ	�x��(��lj�嘻��R<!Q�vQPpcjҘ�1�H�dU*!l�PP0�lZ4��!�D����Uם�]@�v�c�������)Y��ޢ�sZF��[�
;�jtA~p��ό	
�>�?)k&r�9d搑i�31���S����.�Q?�б�����=i��;�]7�}3�7\�)�����q<c�ȳk灂Su��v"��6)y����<�V��&mh�E[(�����#�d �����"�ȵ&�3�E����EX)�f�4!��;N���YJ�mK�O)��j�%m��sٜ��иœ��=�����(�]����]8F#^_�4bf0B��q� �\���)	�a�����R�GQ,c�,�P��/��!e��7m�U�L�P�a�OW�Tu��WmQ�x��fT��"��ᒢ;�BYU�z6c�B�@�_YA !!^�]"�qŚFf{�Dh�9�� K��S�ՠ���p�IdD1!��\?M���M����-��ev���y���+�iJ��4,Y������G������e:�.���Y!N��.R�բ��äڒ)��\D�Bn��ִ*<��e�דҖMl�9Ʃhm^n�c�*�T��ݫIt�j�T�¤i�V�.j���gW[��Cb\Ųq0�U�g>���U>-��~\��9#b��šݖ��]��B@G�mt