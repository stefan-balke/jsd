BZh91AY&SYNzi" �߀Px���������`	>��ysn`   f�u�N���JiA3iOQOL���h�z�� �A��	M	%6�� �    ���a2dɑ��4�# C ��MM42 h4   ��G���&��2  4II�L��Ѩ�24 4������VH�H@��2UIįo�ث� ��heQ/(��$R�4���(��Ek�ք(�h�j�*B�k]������Ǎ��~Eʷ#r�T�]CЋ�Ȍ��jh�܈r����D���\\[�ਸD����7��5m�߶�8���ׂ(����H�)���y��%]�'�\��e�h�����Fy�is��2j�^TI��T�5�2�$ui�Ey��m�Úf�{�F&NU �R�5�³�E�T������f`������W�{���{��t��&�6^��x~�цa	&B�_��8ov/lte���Ӌ{+jf��0�;Z\�e�0�d�K�s��cS�j�۶�1��.^C�è���7���-:Y��J%���;����ԁhg��"�#n�j���*Y�Nt<>X��]�\`nb��ę�w�t��4��3����\���bQ܎�
�WTW7�Y[��ymC���g_Ow�I�X��@��)v��Y5�NukC�ӕ�Y��=�9Hq	ܕ5�6L@�R5�=��m	�:rkZ�X�p�9$ɖ�
�v�C��CkRĕ���Lj�ꐬ)>$)�\��j�P�Y"�Y�L�F��U�Up�Ԑ�8��T��1�,v�VB̈�n�m�6�{x}�B"fU�,���*٩��d�{��xaH���B���*�EJ��|�
���=�������]adAu����挣�9@�y�f4��IxF��1,���e(��~:bb[��|�܏�s�"JӚ� j5�MXY�6�)!����R`5v�~]lU��qFZG.��l!�c��K�䂇x���m��#��Om�V�fl�R��֒���8���,J���nfڟ�y����PR���}� ���8QE�UV���!ѻ��������uN��f�"���:�Px��BH"�H��lPQE
Z1�4J��&��	(�5E#I�Q\	��p6YE�vXX!�n�� �Azn��R�{���.͌��>Xt{~��t���ˣ��������	дDq:�u} ��E�c�������^_Hl�����wwt�T�QS!��U�G�"���u�ZU*N��I�(�P��]������b�.S���8A�[�E�7��
��n�a���9�ф4�P�=E�C�E4-��|11Jp��=���-M�O��K,���I+^%��>w6ȓ:J�TsZ$nw��U�K7�ъ�.{r��H�)*;eD��#�Dդ�Н���C���f�l�UT(j�lb��}~U}ca\4�-��b�2_��Og�OL��#�s�y�^;2�v^�F�R�U[E�ME��0jͅf�D�pۨ'�]L�koD�mSu$�-���4�fYe��ꊍS]I	ӗZ$z��0��e�W�Tn���5:pI�b��I#L�U��/n��ΰ�wn�d\�ec��Z�YjI��1A��G��Ъ�,�؄���$[
QZ���<�"V�w"G���Db)��؄�Ҳ?�6=|�յ������]�'d��wW�t�%1�w�ב"�x�����Ǉ�։L"F�٥���SG�#Q��V�.K�RcHKE�n���$��n,����Zeh˘ӥ��;�a20��m<��FM7R�S��j9�-�'Z9�.g��G����lacb&�*kM��~��5��XU8	o�J ��LP߅4�I/p�c��ET��Ls���c���@�i`s_g�]��BA9餈