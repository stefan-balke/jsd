BZh91AY&SY�5� K_�Px���������P^���.n��������6�h�0������h�%$қ'��     !!���FF�&�C�OHz���A����A�	���dɓ#	�i�F& �"@��)�$�)����j h2S#�^M z$��Y���=����/tA��I�XI�״?�6�z�	dhZ4aG&��������xz���êx��^ŗ�+II�#ߟ������rR�Q761�c/�e��}�QO�n���ar�I&+⅗�"�B���E�H�0FelBi�����	"u���X�KE�B��Na(����֦���$�<�>n!����d]���|�c,�"��(�iN��o��6�9��7z4(ù�:C�z�Ƨ5�AfJ�AEh9F�m�$�T��(��dZ���59�V�I�:�U��,�lŐݢ����,����]ЧY!�6&٩Px@����"2�
��z�p��H���W��|�c���m���Ϝ��]%��#�
I�vQ*Q%�.9	'�K�����6�#d���]�Cҋ4/.2�@�([PP0�p[o�b����߿�;��)�m��@�a�o�W@ެc�ď�����:��Q�����i��*
/4R��@�SP�MIb$������\�~!�ט; ��!@�C�M�����Is�@�����/anFC����%�]��x	y#&f�
	�������;����dx�Q$��%Z��'sKq��^Y�2d"��뎶��(���Mg�K�*�>�u�d83����Y�&�@�9sC4$c �+ e��G����(�1/4�"K�$p�<�k��fL�*����e\�����|�>W�2ÂO��a8�b6$�ؼ�B��tZ���z0X�����xw�8�{G��e@�rp,KDT``L6�-c�1�=�o,�� (��PE�;�X���ЗH�d+��h;X�dF���T&Ȁ��Y�B�q��	��!.�L$oL��?�%aI�� li�q��R���c�	��v�abI'�4q0���%�M)�1Z�s�pv
�3����ci�8Td�2aH�&8Z�~�Ш̺��U�WXi�m4���MI�����J�� �l[�A��iB��$���RX�JUA���U�4�>O~SI�� ���50:R�cl٬�b�z@~�\���-w���C �H[���H�
?F��