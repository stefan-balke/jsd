BZh91AY&SYvQ _�Px����������Py@� �H��i��OMG��M=@�h��s F	�0M`�L$"�&"6��1<�F�6����b�LFCC �#	L@�� Ч���$  =OD� }�H�BD?��:8�>1Z0V��j?�$���д3L"h�TH��Pl�>������c���g�ѭ�xڙD���{�2�sr�%v.�7|Lwj�2��|Y��{s��$2eF���Ȗ��ĸ�,��	��B���A���v�$�J:�@�F�}qnE��_.�/Ci����kF�oB��9����מ�ū�-׹*k��:?�[��KM7L>ƣ�=&q�Ì�F�Jd�48p3��0o�Sz!6�6�(�X�M� |��(2]m�۪���%p�ǭ˅+�Y:B%W��qn	�^�5P@�c��7�lc{�m��
��'?�>�W�G*���T�LS5������l0M"�q���5>vP��kP����ay<ؘ��Z�a��/�뇍t�+�6��v��H)�ھ�8�="�h��0��Ulkf�_F�fJ��v$
����%~v#Ѽ>0L�gI��8����aB����*��D5�9��e6��e�z���"ə�)���J�cl�6/�� y��I:��銝5�Yj �ld#���Ԑ��0�Ġs�v�N
30��K��3ӁY���	��CC��G.a@�a� �Y�j+2(9
!2=�x~���0i�6]dQ�r��pW��D��9Q:������䰢�1U��#����"����H��u�(B,mkh:�2
�t��%��D0�;@T9��Y�� ���
��ܕ��UTd�w�u7!o (��("��<f�D�b�	���Yg0���h��(]Dd��/v�'�M{;e@@���DF#�5�V�q� ��6N�ȱ<*Pk	�f�Z� h�0Î���T{�+
G�V���a�Hm;�3~�$�pDGp���g���8"v�V�D�A�*Qv[�$���@��e��j4$�XV�"����r�D�yv��}�m&�������6"%��b�(���m�;omy�)R�՝��:
��'c'�rE8P�vQ