BZh91AY&SY���� @߀Px����������P^:n���
J)��S�"x�S&�1D� 4@4&��P h      �a4 h4�i�  h � �`�2��H��	����DOi��h hF����!� P	*	D(?/�r3�XФ4���&��6��hJ᤬aQ��Rr"��g��}=r�Ϊp�N�q��xO*�D��@^�����`$�����7n'QZ)%�u���{:��-�	�i����"���������6K;�� �hx:���4�4�Σs��m�sƘQEUEW�E�91+%J�xq�%7O'�&^J��*T��ZQ[ԬH�=o`-=e�{6���"!�S ��P��q�}����#�q2�k�-����PZ�a��$!l���"�@�Y�3w.\9g,1�_䫳U	;"��1anht��((懁Qւ���Bak�����DFG�0�-�Y��i�HBV�I$� q�2g�H�Ð
�����4$��ȫL��\t�zHuTD�U
��(a��D΂ĎMP@@ tڭg9��I�+%�!~�>:��I��ɠL�������D>��!v�!��t�%>_[�M�xե�Eb^352+"��Tvv�iI�����K���9"��������JbVMH�L��4I���`O�HoI{
�I��͇ƁD���ּ�T@�f�A�P��dx�w��T	Ye��,-a���0*�����{TQ��� �u`��N��S����qC���L��B��¡g�? 3��`h-21 ��q�3��n��$�$D��ťjc�������
��lCFiMk�qE�3��	�@��X�<���1�%nKD�~�zjǕ�Y��hḇ�Z6$�9�h�)�?c��� ĨG@P`bL34NfAd7<�y�	+�GNJH&@�Y�DA�(�@�%c6��-��$�R��EC�*����ۑ�jՎ���X���!Qy\hP�9Ru���/e�����x����3��s:B�� 3�E���,���u�V�iipZ&q�[�&�zt�$@1w��!�q�1��y1Vda��!��0�l(�2�L�V�\YL���f�Rkq@�a[�H+Q�ct�8ȱ	��O��`e�{r64��7q-��"��yb3�n��݃k��T�m����R(*��?�ܑN$/�a6@