BZh91AY&SYuNP ,_�Py����������`���;�t�� �@$��Q�OM�<��D44z@I���hSh���       4��)�hLM ���4  		�A��� h42 j42i�# `F&��4� �D�FD��4Ч�c��4@di���$��HE� �  ��j����\� ��M~�śp\�H���4r��&ؑh�����xcӋ�No;����w�32s36�m�N�m������s322li	謙"=��zSꪽ�z
9�1�)���29��w��&b)R�[�m���xtu��|t�tʌ�#X�H�y�����c�GA�Om��rVǩ�bBEmg9�
����/%bY�Mk#��{�v���(Bb`0d$�t0�k�~͊��j�mr%iؘ�Jd��N��hI�N/�R�E$�aiS%P��{79�$�c�SzI{V�Kr��k��M� %3
�U��7V��
�F�� ذV��C=� ��F�[��Y�b�֤���]DB����n�2�ʲ�<O2S2�û*GEPB4�C$���LW�
6�Y��e�aj�%th�%��qP�e5I�!����[S���rƗ��'g�5�=�Ch�F�"3����2	�kT�&
�肶�qu�n�eKM�=R�X��"o-��7jVɡ���1��C�:�%�O{6n��8ڵ�iGb�8���oUEg&���h%����5� �A��mHP�����B��ʅ w�4J�Il��2�5J��q:�TFA�H�G&��M����i�6��M���(�wh]�Xj�@֤B�QA@�5�h�D ��@شjz)��y���0�ߘ���<r��Z.�����FRF[s���¯=���V���]'��U�/��la˒�p�J���`���5D��/�Ԫ����>a�B�����Gq��O0��C�$�xjA=�k�3���$T�_$l6A�|jI��^�$M1���:���� ��x�T'k_L�6�.���A��DP��.Q($p`pL2\D0j�D�hR���uZ�8�����M��cC�e���_(���W��5�*
����ڙO% ЅǍ�ɯ$p�;:���� Έh�SB��,ZMg�AF�#/	?�@LK(�ܶN�-��\�D�|W�0�z�Z�ϵ;�b���r�����%;G�r�΁y��Е�a����aXnx�4�F�ڂ(,A�;��{	C.�p������5;�,��!D��߱ې��f�/҉��F�(G���z�53j�LQ0<������>��hL����,HHZ���@0�9oB�h&s�,v�Ipu��B�!Q�聜:Hc6��k���Q�#-��Pf��
����FGE�X��'P���G�B��DD�Hi�I�����ؐZ�A�7Ij�%*��c�U�>�kI�w�o�.��H��٠��|	�C7�{7����-k���w�h��I����)��r��