BZh91AY&SY1=#  P_�Px���������P^q`
e���#�OѣI��4hhhh� 40&&�	�&L�&	����D"iOMC#5@�@   ���&L�20�&�db``$F�2�z�?T�)�f������MM<��`���IPH,�!��~���_8AV�&%4�$ב�M���hX��"���a��u�F��]M�5�ue�Yk�A��R���`ܷ^3[3���N�B����-2���&��������ʋ��&�U���^����a�Rx�ֹ��U݂6-�|�B��\�*��j���+|��S��-��$�;�����r�[��K�I�3ID����)v��}`���W���s�5�^i	�!���.����36d³���V[,ip1*[YV��QDg����TőX��)�Ih��A"7�c+-Um(�D^�P���,_Q�ö�J�sƾ�r�V$Y��2u���5��3��p�HBZ�I% c9;��w�#��j��IQ
�z&�%M��W�o��W�$�4�6�F�lHdGaCA�@��I	G[Do BH5#�����W͕�jB�1 b�0�����>qE)�p�!��c��<*�>e��|�G0xٿ ���qn0�x�x����D� �N�[�_�?��~!��F��� ��5�O�q3�1P=��\L���6%^+�g:KΚ�ĳ;�^h���ΡA2�ו�i�d3"���!gbI�aP��N݅Z��um55L�P��F��(1s� g@��W�+
U#��Eu!��.%�
�z�m����9��c�����fKLUR�}�p~
�`�]�K�$�j��
���� Ψh������yE�)�����W�0�@�]��(�$��� �e�kp���Z��*toIw���:
􏩰ʁy�6�Z�J���0����B���a1%��a&��$(b������	,�],
�(�h%Ap!ߊ>�T'���.����m;J�Or�:l(+g�-/()��Ј��v���,$ � �&� ���X�ҙ犸��:�C��4q�H&6����2C0�I^�V�Ш̹4�*�+xiz04�E��Rw_�Q%R�&@n5�a�jo(P��I�.%%���U_?SH����9My��.`f����@�H��H56�F�K-�Y�i24(�u�O�]��B@��