BZh91AY&SY)q�) �_�Px���������P��@�2 �OA S       sbh0�2d��`�i���!�HH!C)�6M��4�i�F�� sbh0�2d��`�i���!�*� !���SOSC	4h�h��d�<�����O��~i��|���CH�S_{�h�u�F�B�̰�G��u"���:<[�w��],��9�S(��_�������[�vt�:��U���F��:qw�vԹ+�5��٫%MQ5��;+Ye�ۯd�_j�uO=pD/�,l�"����)���O��w�Lz�����h.Y�6�D�
\�-eݽE=tK{ſ]�Gs[HF�I���t���lT[-\2���ihe3f,�Ղ=�lȭ]�u�M� ce�ѝ0FB���.�kL����f�|�e�s��lcz6�mD!����@y�.�)�P;�5�]Xv�ߘaL�,P�3.6IUM��dil�-P5�֨(F��\ɠm3����ߺv��L��Ē� Po��~#���P� �u���Ǳc��a�]�g��|-��f�{Y�4㛓�k��֭D>��p�뎿y�S�;a��0% ����z�CL�EgY*AmC��uyc�/�1�ڸ{ ��<�>tXX�p��;�W
K�Z���|<�'�p�cMo�� q��_����3".WW�j�ˣƙ�i(yX�_V'k8h]�&��z���=�HL�a4͒�&���:{���Ø�^�+Ev>���<�I��*ͥ%�B�&���3H[�0�jF�E�eo#�dV�+t���_A�ԻL婶�5F�
)�<6�:��뼼w�a�8�Cm� ����0�ПL��a����r�$kVj�W[��7m�ԵrZ�&�PX��,:$#G����p�*�����c�,`<�D)\�B�o����,���t���삤��W��^{�ol���F�����>�D�6����t��ByɆD��ݺb���4`��u�9���E��� �*�&�ɪ�5C^�pX��5��B��8]R�v��Q8c�d��)���5&)��8Y}�/V]zN��k�Y���|��Ɉe�;�:&"Q�Q����`�T��1[�B��(|xe3�|Yu��lԃD��[�?�w$S�	���