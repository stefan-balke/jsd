BZh91AY&SY�9, S߀Px����������`=�k���@˂@�P�Sԛ$��6��р�� jz RQ� ѐ   � ��mQLП�20!� 2 `HDF��f��h�@@���0L@0	�h�h`b`�$Љ����OSF� � �zMK�$��-H�� ���}��]�ֆu��JaS�7��'�` �h[!�0�!��j��A�<<����t��0���|��uPp4p�S�19"D ���[)
���8�~5g�ztH�J,��K`Ҩ�����!1�.�[Q����ʗ�mG��~�`};ّ�w�q�I��GD�B���r"
yE9<��<l�_��}s֛�<�/tC#4O�*4?PCD#=�9qӌc���{�����S�%j}�n�$� ����׿p)T���%��	~&Ly~�o�_�+̓�9���-���i(s�
h�*'�ôX��y�W4�(�4�б��T/��BgP���i�hPC{;*��-\�n���p< �
F��mY�#0��Qs@"7QK{ĉ��o-�T�m[X�����&��j�X̴��8|Kn�p�e� D3N�n��X��YVM:�M�[4c:\C��J�ݦ���v�Ay���!E�X�×K� �M�Y�-V%vW�3S�Ы�&B�0B�3M�&���$eC��f`v���Pr�Qxb.�2�6���lD	��iP��6p�F���5�Gt�����^���Bn.ƛ3��q��֍�"�%���#�lcc�m��BP���~�{�/?��%Z�Г��se\�:vf�4�% �#E�wUl�llE�2��WT�# �	HmE\H�fF�
�E��\�pI�Ch`�7��
�|YK����1�Br��g�ψ`�J���8�{��@��n�5I�_ۂ�f����1���1��UU*�m}������[�E���8֑'�v{�]��x��zRMT�?�б���W��V��ĥ�π�>�����g�$��(��D�1��_�'s$���)����8���zie��J�lqϓN��B���N6�����4���厦����$sk�4���>3e�g�g���6:��i���[k��fe�z�º4�M���cؿ{�>��-ۥ�<�XN�ٔy�r�8���q�*1��8���C���s�^�݅5{�q5�������4j�)$�b�I���Vܲ˿�(��9�H7�Љ>~��T{�y��0������D�C�s]$��i�����[R��4 (��("��<f�D�bK�Ha#I|�ЦJ��/���2$��(��'���bW�'��%�6=[u.�=��z��F�Saa�峓�>!:dm|�W�ਔ˵��3a"J��%GiE��"M��N�.�ә��w4��YuT�hS��L�1�F
�)�-��N���V��� ]V�l^B�=q��N(q���k5*Z�G^Q��KF�D��7&���(�F����}ձʤ�$�����8Ę3q�Y$�0�:z�;�UOD�=�o+�B�*&�w���rE8P��9,