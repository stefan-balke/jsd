BZh91AY&SY*�c D_�Px����������PX^g����Q!�a�="=#@z���� i�� ��*mH4       		��I�F���Ѝ=@z�  D�& �4d40	�10�@B�5�O&��O5OI�@=G�ɘ���D�ň(@��{�WM���&%d&S]'�͸-�HX� f"h��T������g������4�O�q�xcL�m�}n��NE�߉[�yjn��AM5+��¯�k���)!H���L0�q�q1'a9�{�B��A���u� U��$T
ʐK�Z�^�T�+���K(��
�К`Ǘ/�r��γ,�����VLt�"۾���21c��Cыr�lE4s�>gp|�����״��Eh)r�� J�z;�+�r���!p5�eT0�ȭTmP!�0B#C� 4J(�R�Q����V�D�(�h�.�fdS6a&Ap�/(�j��_���D�0N��v{M�61�m��%):÷B٬�T)'y�T�K�;`dP��H���.F��%�+#(mƑ�e^�cJօ���Cb���@��+2HނH�/�܁zP�޹��d	q���:����-9�EWq$jD������ ��G���7�!�E��$0�j[�?��8��tT81����\fW�xH��FF@B���`�Bk�)O�zݢJ�0_R��L�zL&�3`n_�P��3a�yw22ϡ$�F��ٙ'cK�����C�ȉs�-gj�2�v�v�
�!�Ye�����\��[�pgN�yc�!�4�D��P����=v�.7��R��#�}��;��-� к��f�Iq"�����L�v�đ�s�Jh\�}
-%%�H���ku�Iꜭ���������SZ�`ܓ�Bך�i���~��q�l�Zu&%�zA�� ��)
A�c'yJ� �F��PX����%�.�h���nRR�1E���*���9��r�	잴/Q��������}xU���L�q���X���6	��9¤D� 5	��c^q܅�M)>9+K���:X4[�@���s@���Dc$��G(AǞɌ۞���E-.X�V%IP$��4*Dp t��PZ�0Ҋ�jD+Q����&2U@ї�����瑹��x�::͡kA�.�E�k��E4� �t���s��l�Y�h6�ז��H�
[Lc@