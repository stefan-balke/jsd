BZh91AY&SYA)� _�Py���������P> �8*��S��O�I��#j oJ4   Q4i��h @     ���d� 4 �=@   �L�1�2`� 4a�&ɦSI�	��  �5=&
h�	�*$�"����C�UhP��2M|�a8o�b�B�e� =MI��V .}��\r�㣱����+��L����.�Uk��S&O)�c��S1$���������,aq��ay	�d^g42��Fk�Ϡ�ε<]�@
��+�Ә��"P����L�l�9����-��p��	�hR	v}��S�)�f}&�^6ф!�4y��b���d�*�QY��Q/(�d�V0�.�#�b����9�1�@�sS`r��P��I��
�1�*84,I���$�{R��T�a�2��<HBB�$�P("I,�)��#�P�,����.Y3KT'�TI�P�%
���-&���C�$�E�19n$��0A*5n# D	BA����ҳ�xk��WV3����*����)�(���!^�P	L�o4v��O]��׶dj�V��,oAT��_>iQX�Y��T8i�f4�����6�A�!9�љ��P=��*VL���Z��e�I/*���0l<j���`k_P��f����2;�2I<��l�m��L�v�/-jL�P�;㩪	�A�3{��D���JH�ȃ��&(��T��f�!�N4:�F�苘
�q;`T��y1%�ux�5I��A����#���ξзV���h��A �а�,
C)!�w���
�+��-m(�ykǢ���v�4b���Uw��>p8����j�f9|K	u"�"a�Js4a����D�� @H�@��+"�_�(�@��6��s�B�&����M�mк��'�qn�^s����Б!�����Zf3�LB ������ǜ�H}��hL�#��B�� b��� a���
���pή,<ǜ�;n��A�9�f��$1���"c�"����kۿ!V[�~e��d�	�&�����*��73A �jn*�B�ZH,�b�RX¢>�}�#�݉����A˙�.`k�K1T��m��n���m[
�w�q��
�>�.��]��BA��8