BZh91AY&SY�{�4 8_�Py���������`>��`�/o �!PԦ��4d�M�b�jz#L�@       2d�b`ɂd ф``��SeM bh�  4 ��EOSa��OMM=G�M��6�d�@����2b?E=2jd�M  )�=E҄XyY*%(�7}��@$~]�H3H_�	Ti) �	�\��m�^S@�ƒ�e�B�t��HV������9�Z'H鑕d��{�P�Yoj
@P����7�7�U��0�h�!	G�6�̐+��;O���ݶEU�YA��X�y�=ㅖDG9�XO���z&����'0 ������l^�^W8��Ay��KQ�P14�ǆ���>�E���r��#5��vQ��QQMғ���*G�Jޢ���W�9��J�0H�fpƋ�Zaz��A�V��*�	dT���&RЯVEb�]d֊����t8��=��Ӭ������N$�6fi"#U��6IN�&�̨�\U6I2�"�`g0�B]BP�X
��0\0�J��@mP�)w5�[U� �"�B����/
��Z��ְ�T�3���E�VƮmz*�ӥ�5;�w��cٓm��4
;��Gh��5o�L��K���A�� �E����t�2%�V�"���I���AFUp��E��^P�@@�t�f� Ɓ�hk�4I�_�<n�yu�ó�����']��	����AP��CDI����H
�]c��-J��ӏ����j�ܴ�F�힠:���H��s	(�_��!`Y�?������ �2RA�Dl�@l$�yU nx]	��mf@�N� Gh�� ��4��!�Z��0�k*/��� �,v�4	V�.�Ui��qXjf���E	p0 �0�&P�s&��Α0a�y"��;%��i��g������ ���2�.��W�<{�4=��E�0��&P��x��)�i�����R��*�Ox���[	���K`�vm(��A3�L�����ڍ=�횱8�\�b�4(ҽv��Z���ԚX��k����=�:
�C:�e��Ȳ��D����C�V��d�2i�	]��aP,b�N���*+�<P��Ukp2Ü¤�EC�TB�� %s��V�9�X�����!@0Tk�d	�}��^1�F@�4z��̯:L�8VB�S��fD�c:����0@�P
g�j���u���*-!A�恮^Q��0+�i�A�*3f����"����"ą"eB��`rX��Ɖ�!�E�A�� �P<NJ�鼒.�`�JH�
�@W�,�op����`]��]c� �e�a�T,ͅ���|�j�y�B���ff�150��§U���H�
�{��