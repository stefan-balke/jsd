BZh91AY&SY.��� �߀Px����������P���u�6�Z�$���J~���OS�S���~��jF�=M4=A���mJ        *���
�hz�P ��0L@0	�h�h`ba"@�ML�!24 4  4hȲ�(B�.��J7?�thH?qI�R`�e���śp\���@h��R��0�1}��_�[��mu[Hΐ����V!��d��g��	c�dJP�1�'=#,�sZ�.����U��2�,\b;h�dC�5ɺZ%�h�͈4-o;��	B�'�
`�,��u�fOOOS����q�#��L��0cϗ���GY-�9Źm���N��C�U*�ra��%dn��&��ۉ^�_4≮ˡ�)���Tf�4��!�1�������&�R��&�P�� ���(��Iങ �P	5�qU�]�(b�5���I&�`ֺ���:1��f	J��M�؊����l�!)B��e
����3��7�lcy�m���B�76j��a�RN�R�-v��L���1դo
��t�J$i���H�d�@Ƃ�E�u���2@�,~����uO/��j�kqa�� ^n�����o HS$���L�������)���ۨ�Nıŷ^�c�@�-F����oK�4�/�j�)��� ���t�=�;���R���N�j��@�8�XҒ:W��s$� `��D�y���Rf���d)����O��A"��I�J��%A���;7�7hPid"(r�-�Q&P���Р��_�0�l	�g�ΌL+��6��˛�P�%�7����Q-�"�8%��6�B�88ƉrJ��2k��\vG7-|!�F�2�!�K�B����
�H�EI@1��v�?��t`j]�i`@8�]z���Z�6�Hb�f�%z ������y���pFA�+&#h�03��+�<��� ��{Z�(V D�`{��\1U�
���R��EC�XH���˳��Bl��q� �E �p�^�'�U!�_�a�C�̯�ã����q>�i�'$�q���I�(0a��lh	�3�B�X�;E��+��2`N��x�g:;�-����lo*3^��������H�:�ԞK��*_!�C6Q���P8�]�Ă�]��,s�y��F>e]�#�ى��h:7n5F��)8f�ʁ�H�n�FۛG�֩k]�f#A�`Я���.�p� ]3_~