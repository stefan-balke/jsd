BZh91AY&SY�r _�Px���������Pf�Fx �ԍSz#I��4�h=@=OS@ @��<�dԁ��L� h�BBL�m@dzL�@  �h`LM&L�LM2100	&���# �R=5�=@A��6�$��B".�2B ���|GA<A��I���S_��ٷ��,ƅ�fL ��j�9H��{���f�׆�������D��}n6L-O<�`�Ƶ��H�5�
�d�V�qE��:'e2�L���s8�g�1m���Fq� �5a&=�E6D�9=���xeL�
�zr�ֹ��R�] �R�״���gTn^�-�IҮ5�3�o�z,� �0��x/�di�2YT��8�W�Wi��yy̠8Z(xm���&���6�f3O-o;eg)��ch-��*�*TߡmVUc�Ҥ�1�$!!	M&�hi�	��*K�� �B��<J�Ir��@���ܑ��,[""�*A��H�2����(��aӁm�i�!�ίȗ�;����/a��M�R�>�5�8�jc�� ��Q1�h��n�쇿{�}Sپ��۴��$��i2>���>k���y�AY�1 ��{�5ݬS d �@+��eֿ���Iz{K�M���Y���	�X��hSD32���Y�_4���)]��ƌ��u��͐��v[7RؘphPu��5lUE
T,%��5܇>=���GH�8Ĩ��+
s� ���5���]�������dIw�G
#��=�f[��eD6$�4V�kՅ)i)��������AP�U��ؠ #J��.��:tݵ�Hʛ�yt>@8����ʠ��p+%�(00&�1�f��7<g(��q @H�@�wı!!���E�0�3�3!�Ċ�@�d@Ee�q>U�	�V��`3�<H�?+���^6��y�C�cBe\��VI!��z9q�F!4L��h+;�a`r��!P�s@�Hc
�"C�Qv��Pf[7�!�7�^o�Ed�Rz-�T"����f%���5�L-�����7
�;Nғ�0�Z��)siz�XM���a�h`f���J	"��>�mf�Uv~l��B�
�Κ�]��BB0@	�