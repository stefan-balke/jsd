BZh91AY&SY���� �߀Px����������P�rB�`A@J�I��F���4  �  � �`�2��Jd����h�������� 4�`�1 �&	�!��L���#
`M��S��=&� `M$П��Q$��@�����`�� �LC_�6��1"�\2� hڢdm@l0[3�f��-�]B�v�H�s��V��|6)R���U@�՚?����V�Q�.1��:H.O��]gY���6�y�j����4��_�ԢX.J��l��xYt��-��7 �S�\^FyܧR*V���I	75���r��w_x�{2E���V�߼��G:	X]��cL�����'+}AdDd��(�ɕ/E���bP���'et�R��|�h����H$N��*K��;�0&˪�Sq�HBB�$�P(3mN�0k�7s9d���#�#u��hj%��LأE�� ��uP��r!�.K���@�k���!@��,�/���w��ٱ�g6��-)�c�j��PA&�gg��{�mx�0d����%RY1WW�l����5��B�P��AQ)M�(4�<�؋�F�� �u>�׳b�nBܼ���s��͜i)��>�>�ɛ��3sZ�Y"c�k>�_k ��]֒yP%Z�}��?��Pkd"(t_.PC�4pbPK�C�E+
U&KŜ�҇>=�U��bq�C�XX+���}���/3TIu���;��ꞥ ������MuG-���^���H���T4a:!nuۼ������������-�<`]�jh�p̏���<�Z�b�X��-�x���4r���]�10.%�8������Cs�oI#I 0�_2	
U�#cPr�u�*���`nsS�AI���XDM���V�'��P'!0��̑	]�7�#j�7|6���r���A��XЙns��@���0�vm �L���\\t����E�i�@�NA��S��1�2F{�Q�7[x��`13-%�\�Xc����6q��LC���@�u�$�å�K<�S,��?�S��g��fmi1z�8��{A�:	�����H���Æ���AKZ��CA�`д`]���"�(Hs�D[�