BZh91AY&SY�<t� �_�Px����������P�n7`�@[%hdi51�6���d 4 �Oʍ�4C@ L�  	OQ)�E<Pz��5Pl�� ��@��b�LFCC �#	 �������P�!�G���	��i�$Q Y������i��0EAb�:���9�`0E�^����&X�����q㧊�t�K���W뤢_�H�ź0t`ږ�j���?y$������PeK��Α��'��KQ.������A�b�<&��k�s�T,��2������Lg.i��Eݛ�a�C�c�%���'�ay�A�	�'G�\(�/�}M4��jdR��ՆQ'��IG�� ������C:��)���APղ
�I�*���a\z�!#�����e�wڒD�p�H`˫��Z�FL�\.�&�SDQ:��1�o���8��^B[��Q`n��X�M��5vAVA�z��dn��־�-�a�B�A�b�%2Z�((�8�Q�P̜���#e�5��Z1��g^�Z��4ǹ��������h�
*�k�"L���vC�je�,�paRL���pfq�ػ=�y�;��1�B���ܴ��v�I��/=!=��f��]� �|��7�T
$�FK��66�C7:���� ��w$���[��#���ӆ�٨72:p�mPAf��I2\D0k]|ů'bl�_����e5Fd�ª���҆���^����>K�7���A@T�i����M�ؠ�~z1�]D����诠2̑���*d�$�	�XF&q��R�`l&�S̄]�mh�p�G�p`<kZ��4-+Ua$l�#ǰ���OH���2�^s���Q0��9��a���I�� $sb�D�d���D���$P/	U�
���R��EC�,
'����w�Bym�!�d�f�R	����=���J >dr�!�Ͼ��7	���0X�C� р(��*ڑ��f�|L%DÚ1�J�Ӫ�	���\3�a5�[P����;H�:�ԝ�sS	���iP)5�P3�u�$�á�I��ֹ@я�S��c��boi1x�r���cz��5�r��yt6�KZ�՘�㬀������H�
��� 