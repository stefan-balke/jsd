BZh91AY&SY�} ߀Px����������`�g{z�`��@S��	$��5Q4��ɐh @d�@� �@  C L�4ЄSС�4 ڃ��  !�&��@   ��L�1�2`� 4a����=S����2z�0�dm,� (	�HFD ���������0Ш`���e5�>�ۂ�$���a���T�@f@���Ç�����~������8s
�.&f{�gi�[Rw��o`�x���߀�T
������qF�8/CA�f5��R�H��Y�@�ai�]�^�F����gt��?��s? ������@�6�`8Ɏ��`�HN��"�C���ל�`�jz�$!R�%! P*�CH܅�DN}$RI$'s�T���qFL��CG���L�9l�=`7�;%f�8�7톨@�x��z	��zC}������9�����a�}���4�4��0���U)+�2i��[�t�l��KĎ1	��[F����3�t!��"��)4Ӧ[/,ܲ�zŵb�hL��b�����fB�#H���ΣQ���SW�0Y�-Y���ņ@�([;�*��(0�	���G�!�`�g�����2]ޑb�uf�A�w!qݮ��2*h��eĬ��kI!��
�+�H�/
VG:�0O)�)��(�v�%��
Ί�5�W3l�X[�@T�(�$�웷VZ���
�ma��#	R�:�:��ճ⒰�g������7��Y�6�6�<��v%��6��&����h:~�H
�x�)��H��#�ԛ�̀�]���D$�+m���ೕ���G��(�!�pbʹf�:e�u��n(H8DƛlWF]e���ԍ���tCK�R���EEH2���e�F4H!y����k����lBL��X�t�3h�vY��>�;�9BP����U���IlV1���B�~�]&>��*�'�X��Y=�'��ܜ���� LDĖi��d���qǴr�aĚM|�Je�b��� y�wE��z���5��I{��8*	�-��1.	�p�H��gZhB%��1�.
�#*I/�A�g�a4������$�A��*��� E�	'|�4���Q�6����3uj,�!3����ІLH7�7�$�"5v�4�Y6X?��@�e�p�y�*�x�1	����	8bL��
x���n��X`�(��=��g��P�K��fLd�yq�;;��[��2�3FHY>��{J-�z��=$� �4��S�>6�.���u�k�DB�Р�k�f�1hW� �iؒK��<@h�O���`M`;�A������"���C%#HV7|kz�$�p�@���� �͎�ďY;�0�yg4�ݢ�h*h�T� !&0zpH,:�Bx�MX���pH&*�2F�{�xT!�`61H^/�W�:�|��2��S�T� ;�@^ hk0@a��$�HD��
ҧ3��9�afp��w g"1���a"C�Ё_���f��H"�����RT	(�n�M$�����p�5E���}
�R!Z��7<�_|��a�	CJ��ti�[I��Aq�Z�kB"T֮($P�H��(�궽��:��ј#�vr��]��B@��,