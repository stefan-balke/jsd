BZh91AY&SYC�� ߀Py����������P��e�H`�������Q�4 �    	@�dd  �    �!�ze��=@4  #@sL��Lф�hшd�� A"I��11?RxI��C�z��x�9\�OZBQ	"�� ��r�Ft��Y�P0E�)��6�@r\2�
��0�ړ�DT�Ϯӆ�w��s{Q�W�{q���c�5��N>�����vY^A*ѽ.��m��t䶚�J�f)�q�l��򷿬?Y�AB�\�7Z�.�[w6��}ۖ��)��W4,�U@�)v�Ә��,B�PtP��LscUU��^.?��(�q`��M0c˟ν �P��6&�~'L�!\�N
t��͒'������lT)��o�U+l���|# ���ɆkB<L�7��Y�k(�NZ�֙Yn����y0Z"���}<@�"�Xl�<&�s1�|�X�%���L#�S#��U(!7j��B��^^oj��&�,-� ��\/w,�J6��*½�F,��,�^ �ޜJ�g��@��e��S���g"�5��8M�TQX���m!B�/톪��G*��(��Vcr�Tl��%��&(�yR&�#��].H�2Fl�aAA@�5�����1}�A���Z�t����h |.701��O`juG���[����.��f�W���5b�VH���m���5j="�".�H�iH^`�5o����<c�;D���� ��4�Gqߎ���� �=��:Yz�f[�]�&��b�.fG�a4�����Q"��C0<��l�yg4��a*�4��Xе�z��B0*����Ր�x.ĸZ+X�c/�U`d�3e�C�9v��.�6�m�Ї/&1
0��-�lB����AB\�Xw~��V� �.<flc*]��u����� &cZ4U4,_l�v����T����3G��CO�S���+4+ؔ�|W��wW]z��ZV��H/�B��;@h�O�}nPL3 j(Fԉ�EA�eR.
��S�I3��("���.�z��VH�d�Sx���	XGT$;�#B��z[P�:�LD.��	��Aqh�������9q�Z���6�����	���P�B�G-Bh�a���!P$T��+�b�Q�XE�af���y�3v��9��9)"c�(Z
��Pf[w�*��i��
r�IG\g�XA$ˌʬ����I���}afj
Ph]M�Z�^TQ�0���.M"�7��CI�;�7t��f�$)2Y�ĭ� �������T�K≠h0*	�����H�
q# 