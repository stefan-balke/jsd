BZh91AY&SY�� �_�Px����������`
@Jb �P�zj�'�6��24Mi� h� ��I�T O(  �  s F	�0M`�Ls F	�0M`�Ls F	�0M`�L$D�4�56��MG����A�dj(�C␂�@Ѕ���9��G�,Ф"��um���,F�pe�B;ڗ* H�@b�<�GC�����F�n�r�֙ꞷ�F��Z0��'`�K$�ڇK����M��X۝�k��Љ'Jئ�k�0�	�A��'�|���<(Xe�6���� �<̥l�a,Ɲ�3Z=OU _($+� <�D���(>�_�O�'��]yD!�x���=>�:�e��z!�Pcxh�2	�2`S'����� �a)uc_Q��Z��D37[�֊��T�Y��@���ҪMM��.�F8 y�9Ё���
p��'��sQ!�>
d"kg�Y@ظ'b`2�9k�ҵ�}e�e`�.n�6�p����jb5@�X�#/r��0��b�݇ jmcU�����!'�X�XU���3�U�bM;!���'
t�h7a
�.͛
�n����7H���\^�酵ga�vh���ik/�i@/&Ӵ�3�,7jE��L\[��8��lc{m���� �P��y���bhQ�y�Bi!
`%�4��DC�.n���]����* ��@AZk(5I��Q0�! �����J��������WWSf{����[0�	C�	ף�͸�N�i��?�#�/�r�A��n�>VG#Ԙ��|xrrJўFaS|ݠc�C�P�X��A��:��<��>1�8�z�!�B3��g��=�y����@<W��+ھ9y�Y"�#�!lf��P�L��ܽ�TLC!�������=��'��6��Ѱv0�����`����z��U@ʜZA�1 �������6Q���ڐ�g��\ֱg��H�N4*�7��@��6���`h�(
��zC���@1���+|���J9�B��d
v�Ld\��D��H�(�VJ�	x�99G����~�Sj�.�P����-���=���spC����'8sG��x �B�����n�bu���s%Q���f�R��hn�(�%Y(N�����9"b=�AT��!K3�h�,TR�`���DQ��h�7'�"܂�qE@eL�J�"My�)�A	 ����4 m��}��hL�Q�:�!�F@��w�(���E�s��0�a�`�0��u@�~#$c�"Q�6��8���b�"�����\���^9s��H�!���P�
Z�T6�a���h;��6l�����#�U�i�C���>�n�Pb�r���*Ȱ���9��z��6�ǑV�����p��e���.�p�!�64