BZh91AY&SY�<Z �߀Px���������`�ը�6W   *�	�2h� �h   53@D�d414  �h �A�ɓ&F�L�LL���� �     `LM&L�LM2100	A�`#@��e=CC@�i�2�uC�!@X /(?/��rg����
F�Q-}��B�i+0�	����������r�ǘǍ:]�iƾ��m��2�6�u����+���	z(^ٞ2؈�F�n\ӂ�LI��R+6���^���콅
Y0���F��&�� ��$X�����5�⭄'��MI%A�t^v�
����D�E�4d�D%p^q5��[��)ww���
�W���4�X�mރ��F
�0�xN�[m��
����^VP����_�T/�8��Q{V2¯Aq/�Lm�M�#��"e�+�(;��L�aHB���kP@���"��V�� .�-�X�0�3��=0xp� *��ih]`�%�2�`�c'+�P�P;.�*�Tk"�c*�#M�Q��F�J����8�]��T�4.�����LÜ4FtH�de�2�<�I7��JN#%*��ă��A�{W�b%��r�"�HKd8��tݢ�2D-3�n	��a� �D���8B6�6
�R"��e�\�SuȻ�3A �A�$�Z�Ao�j��Kð��:ǮH���3Z�pӐ i�4�v��R�YI& �zhB��c�.����]L���$D��	�I��`�!!!P�n	���Ӊ��u�o��
���z��
	�.��Ny�ɶ�6����nQ;�Y%�--�=��Ӄ+4&��R���$���w�@ B>��ɯ�v~�G�;RW�?���S���<�b�w�!y�2�i�_��Y~䗟���<���g֡Q3kZ�\Q4�C5��A�]֒y�k]~*��.3�!�]
,�T������2�[ؗ*i	�P��)��s[*�t��6���m �AUɤ.u�� �a�8��QHX����4&8p�j(��G%���x_�qB�!��D-O�Vҫ`gT9��(3/�:�7ԻOsR_�ii(�i�A赭ɷb3,�H\vځ����l4�2�q����V�f��hn��c�%�@r�P"B����!��2*�P�&��2�҅�",Œc�f����GI�G�P ��� ����ǻ �ɰΈ��|�g�mbr_�>��4&]�u�q"��	��f�ց�T<�.C!y�}�Q_�`�0Xm:�f���.QA��38;cqp�[/�+B-�7d��t��QK�&�c$���̳Q�A��n�����9Y�h�� ��&�h�S��1�{15����sH`�j��U��KDwI!����ګ}��4��B�1�}�w$S�	��u�