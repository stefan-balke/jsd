BZh91AY&SY��� �߀Py���������`=�%���@���'�i��� �   S�#))� i�     2dɈ��	�����$$��M�6S5��144�i�48ɓ&# &L �# C T� &�6�&�&j{Rd �jjyM�EwD�$�D��"�W���v�O���D�TF)z�I�Ug�&��`L�F�UAH�� j���l����xy+|��;]�ڻWi�;6�/�	�1ߙ�7����1C� ��f�yq��d�Y��|���q��U����d�M.
¶�Իd��v��Z�9㵻j6�����٧Q&fm��(���c_
���z���^��?'y
UT�k��;�u�I�^�釻�<� yR�J�2D���p]��	:1 }�"��{` ��*���"�M�ق���'���1�m��UH�B�^���� p�H����*�	�Zh�2�0I�{�¡C-����C&�-.!�2 ;�*f�e#"�
��$���6p4V3x��jY��>��#!��A��4�e-gm]�Ų&����k,��L��W"^�<<(B�uj�Zmn�1n�!�'�P��4t������ZÉ�$�6�L�Q��4����o��m�4 �=��Ii�G*$�M�%J$��T)�(1�q� a��"m6aǁ��TY��M�jJ*6D��A�TZa��˔Z�|׾ȕR�U��{���3�R]�]b� @�>W���`00q	�2C�b��P����zx�I Ԙ�-X�A��nA����o)��B��� ��ϙ_�V��	&�*!�B��[�_s��)���iK�u���M�:��S>�'��2$���
s|�1Jt��y^g��'G���Y�h�I+v%��F��Jh���^�5Y�Y�KFXw�eL�Sp�;��d`T�lr��E����*�yw�m�}�E$�pbjwr4���x��髙ť�`�1_��?���p�2X�>R�թXGvq��g��yv0X�Tc|"r��N&��x�y�l�o��m�4uq��Cͫl�RK-�|����,����f�r˰����S/�_eQ�S'y��oiaڍ
��I�&V�Ë�8[c	���Fk�B,;^X���%�L��.�l3(�A���"4\4�	fH�e���J�Ǒ[�0����]H�_&׍��Ss�ia��~`��Q���N
�J�L����f�CR���TS�YF�gY�w1~&��/K��]4;r1l2UJ�����-x�_5����ݬ����ܙZ2�v�ݹݛ�%�N��$2j��c�d�kT�:1;q4iй�jI�����y|�c��2�#wҺ�9Ԕ��G{���RK�uaML���t����U>.��h�ިrQQ4�{4���ܑN$0`y�