BZh91AY&SYk�� C߀Pxg����������P^㻸r;Q�BIS�O&iS�z��mMOP�6���i���OI�m4Jd�4   h   ��BT~T���F���=�@ �=@dɦ�L����0Fh� 	 &OD�=MF� #OQ��@�$��Y����FD��A��I�XI��x~�m��%�в��>6��H́���y=��x���h���&�-�L�/�����{�J�u��6��KK�VT��h��>���a��-�����Rl��4.��GZ	+�ք�Q]$ U
����-#Mv`3R!���ꞩ6[��`��m뜃����r�\ӵ��tܱK�"�x�T��e��[����fi�ƷhC
���3:�=�h;�ጻ����mnƳ�kQq��,�K���QK�PkcW��[��-hD%�J5M"Y2�-U�3�*+��QAq6٥�ZV�"ͭZ�6��3�61���CIB�=���y������e�d�����.�u|��/-H�puQ��Ɗ��CV�҅��A@�5�n~&1�6��|�M�zgѦ>sL����j���y�Q���	��,|'����2��MA]�U�NΨ�����u�����{�b���:K���rYp��)�K���hTs��߅w�!�0��0�b�ZP��~�'ʒ�QH���+4��gB�	��g7�<���;�:�Mo�V1��8'�K�r��<�""��ڼm]&\u1x�+�C���U�;YӍ�pg���z�M��i8��E�@GP��Z�l�JpD~�������̠�ݴ*�Mn$���N�|A�Y"�!�����;+�Am w�N6`
3ʲ�-�,� ����V�ɫJ�������K��� Ѳ��(�9@g�T�e�֊d�s2�a���I	`P��T�X��l:$#�2]"�V�|�hn�T�AI��b�6DaՕw�!<���8� b°\�H�m!��j�8;L��\�(p	��9˂ĒOhр�i��%�&���U��)��b��P��*6�3�]q8Ɨ;����d]qqQ�xn�*�+|.���ZE��&����PJ�	���b#P)5�P.��~Ă�]��,x䪂P�-��2D��2&�2�Ə	�fdI����$�5��k���8U-k�,��� �0d*�9?��H�
u��