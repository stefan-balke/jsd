BZh91AY&SYB]�� �_�Px����������P��c�Î� 	D*mO'�MD�@ M4�	���h��`&�`$"������d��  <�0`��`ѐ��&��D���d��@D�OM5?TyOH 4i��jj-zЅd��	%f�x���,5���k��[ne�ƅPeX@4w5)CV -}[�n�>-�N���u�j�P^�S(�7������+l�kEU$Su�s�\�a��[�C��q0���;"�H.OI�#I�E�b�,]�{iZ�s%Z��`�@��h0���������R>���CL������a���E��8�_d���e���G��\���!��u��� �E|LU�EF.&HC$�j�/.+G�h)���_Q	ͫ8Z���!���zV��ŝ�6��J�C�1�"R֘��1�G�A�CU� 'B��"�"�![1kU\�DHA��׃z���郑y�@tY�	���T�nCX���7��m�4"�w�:�.N�
�E��8�e\�"�7��UT�M��BɈ�K�
#"p�Bd��ui�A��<�/#[�����if�;Uteg4f�#
nn�@� <���o/je{�h����kڲ�2�TD��M �zl><&H���nZ��
��cUl�c�S�M��:B���n`�f`�8�=� 1����3�X���A |��O>���͜TEC=���2f�مb����Z��H�cP�gʁ��dy�=i'��*SE��Zο���Pf�DXt�.X�,�1�+|C�̱`'��|jC�9xM�͝�46�li2,:¡N���=��"VI#Ba������:H�PC'��(91�F5GOE9{�؆��4,߯=��hiSY�?���!U�2�B3�JX��Fax�V�ǥ-�PŊ��@�<{N�9�:ǃ���``T�Ȱ`i&09�!�1���@\�9( �a!ҹ����$��0�3x��ڼ
�(��60|�ݩw�By��qS��AE	��/�ؾr�H~Pu���ǾC�Ƅ�gI�sI!���z�����iL�d�*v���^']�B�!Q�恜��$1�C�Q���2KV��Tf��4���\.W�+"��\	���T�C �n4�C���\J�>���Ij4���V�#�!}j��"��v&֓H��$p�L-h3JEL�� �H�~�l�׶�ͪ�4W�eL�A�`Ю���rE8P�B]��