BZh91AY&SYzi�� e߀Px����������Px�b%e�r��!)��i�P@4h   Ji�ޤ���@    4������� �ďHhm   � � �`�2��*������M�z������@��54B���WI)
����7��� ��D�V dk�}�ۡs�Ig)���4q5"����j�;��6j�^R��c0].7:q���,?��Ď)l�rl�x���j��6X���x���-��r�nb䈢Ƣ�>�Jʢ��*HqQVGR�n0Rժ�3���!@}Y�òiهu�KW�i��o��w�.�1�kmV��uk�M�1�H����NB��_�K"��!s�xti+DdO2q��Z6�-���E�Qz�1�r��g)�6�J5g8���*�X%�F���_DcL���ҡ��ә�K�(|hNFJ�t��{���<��i���c��>��,�4��mƱ���o&�m��(��sg|<P[��x��\xX��#�w�t�U��M��k��;��i�eBPg����)�ކcB3$#�����;�$�)#�%g~`�Dm�����wf8��8���Q�ԘZBkϏZ4b�g��:X�)T5u�X�-ʍ�����ǩ�\��������H(k4;�-H��J�j��G���l�_�">�z!���k�ij%�F��o�X��%�i��TQ�������Q�@��uu�;9��c�ZN���� e�u���D���|)L2'��������
ZTm�I$�0�Y���>o�k'fm��W��T�_C�~���ٌP��Xd�x+ˡ���w,S+�0��B2���f26�)h[9���?�W�쮂����)�.�Bv]u�k�Ǆ&��F������%�	�5���;����\��\��0Yc�Lٮ����(U݌Q
�Q7�q��xf 2�p��^�b��Z��T���t����;�,��i�U({k���knj(<;}uu�GHo3Z��ژD��;�KՁ=�0�%&�{�a`��̽����9\i-L���;�Sl�Nq�u8-K.�Qu!vc�xjp���MőY͟�h\�X����hLQS�.�>eK�H䶹���V�(X�1�S�1~S��b%ܝF2^��f]���~;�st[~�slR�0�s�"��]��BA�6p