BZh91AY&SY�U �߀px����������P�{a�AΖ��͚�p�DOژO$�=@h���ҍ h4�43Pj1'��~�4A��4i� #		L�	�i���I���@ h�8ɓ&# &L �# C � ���LOSji���h�� M7WHL�$��4@@�}����?��
��,$2��͛p]�� ̰�4z�Q� Y�5}\OG/O-�K���0�O���3��5�2����[��taj��"�dܘۖ��uŕH�DuY��m�EFRV\4͢ �As�8�9���lcq�nAz��{�BK;�8^�%��G�:�lk��F��
�g���5/�+�Hcm1���a����do��볍�c�b>-�Ic*���u{��U<��[�؍1�Ћa�lWZ9v|�� 7h��Q�1M��Rs!�� +Q�=/1�Ca�njC]2И*��];�EЊ	�0n#G=8	�6z�|"�DD��C@B"� �d艑L�=�X��Vi�2ܞ[i��ȵw,�ُ|*�e7�uvF�61��m���!M�@x(]�r9P��y�T����1m{ie��	{`�b���!#�S�l��:�CV*��-�((F�;3��0Ch���{v�;:���Sosf�\�s`�M��}��/�Y�Bɣ���?�����4���8}gT�<k�۸l*br���s=B\�$��3�G�-5�̹�C���\�	@�B�cz�N�%#ɐL�ĉ��_ш�ڔ�G0�؋��u�@�LŁ����i�!�ʇ�k ���̒|�
�4���hf�#�uwvo-C�ȉC��d�A-I��B�Z�0j�b�)��+�Ν9��w���\<���m�9�';�
B�F�A���H0+"`��N`���<�$l�C2k��/��:�:��d�P�D�:-��9,��2�&;�Ŝm�!�)��$$k�
,	��һb}Qn�$�Я�$|D��c�GNA�@h�Zv�i��i<�X00&�L����0��I7H
:;���|�tHF�%�.�a��0n�V�qSF�2�d�6;��y�!6��9iL 8d�>�=A촒̈�g�F&�Ηo6�|��hL�a�5���C�����f;���D�������:�f<��Ӻq�Q�����fdTf�r�*�+per[�ђ�*z��0p����77����E*���H,�i��,���؂��.ޟ��.���I�d���^"![ �C�IL��A_$A�~�V�k�p*Yf�ɘ��B�p��w$S�	
�Pa 