BZh91AY&SYwO�� ]_�Px���������P^�C�s�@T�S�H��C@�@    i4�I 2     D"Pi���� =M  @`LM&L�LM2100I )���L���� �h�)�5���pKI$�He"Y
�>�W:C�.Х4� 2Z���ہtP��i+������a=|&���kV��/h������$�~����T]d���YNXۓrM�,,��W.��˖w�S%�~6�гT����ؾÕ���ވ�n���|����Ș��5Џ�!5�m�ni��,�`ǣ�٬9v�2X��bt��,>G��%T�5J�bк$�*�em��2hى�x�q�ZA�Ґt��7�u��Rk';ӋN�W/4��7����X�)��
C#H8!�V��X,]U������)FB��L�đ`)̢�@����׶�k�E���ln֔O�g�C�m��C@A��j��R��C�4����z&��拵q��m6ٸ����J���L�I2ZR62FT�e(��$��k^l�bcHl3gLg-�}QˋX��J��C��!ߟ�E5�%~{�&ɡ��/�;ne��<}��)s���Q�06��g����?��o/9����o�zC>j
��o����{��KCK��>����S.�'�����oo��呐�]�딾R)jqob{�)e��?l��`]�9�n��UgC��{[*�r���:��SLuҤ)ދʟy��r��%�o�g�ZEYO��f�5S֥UUUR�U��w���̽U�m+����ͺ^�0]�����a�l���q�t�]�Ǘ�>�|:׬�Tau�8W��&�����
j�i����3�G�դ�P�b�/|�*ߖX��늓d�Q'y���{�G�����05<�.�&*�T/����W��l)$� 	8��!D׊"�iY!�A7g\f�.R!���. �e�[_V��:�W7���/����#�wݑ��rt��m�^��y�W�nTJa��s2]v�GyJ)���6��=�S7���w�~�*�_
vv)r�&h�V�5�ۛ8�o�Lm�9���K�־ڵ����Zʵ84�*��Z���f��5ii�(�t�w�_��l�WV�*���Y��p:(q2q���m�g_;�=uS��e��M��⢢j�������"�(H;��� 