BZh91AY&SY�Ť� �߀Px���������P��:�g�b ���A�P��d��h   �6І�  4  ��  ! �I����yO�=&��z��  ������&L�20�&�db``
������*{&"bb��4ښh dh2)���$K�B�F �
�|5Y��a�P�BMy͛p^6H�B�fXD�;���D��c���7������M1;�c�2V���L�x�~�]L����H����j�a�O[�R������|�Aͮ����4 ,�g�b�[�����Ө�I,�E�\�L���$%����ą����;?��DB:75���8�g��0dAE�:2��$�>�,�=.^�ќ&/S���o�*A[�%`};u�ZM���<P2�J;�Y��&�Qr����K��#�ެ��)�\[f�r��{�#	S1gH"� @Q-�4Ԣ��ZK
5a�5q���4j�1�B\2��CZ�k2�g��RQ���@�p��P�yL(4adV�Lm���P<����k����3k\{3�B�F,w�#c���m�����:�A��]��9P���D�D���ӡ����4���+%Y�Hܑ�� 6���Ue%l����k���l�կd�M��T���߯��ݸ%������)��u[{ r�XR|S ���*�=���)տ*�rI$Q�q�b4��3�ܲ��$}���n3���}�|���Dи���Sf�T�z�]�l���ZQ���|��$�=�c	��Zs?��қ�n�ݦ0L�����d!�g�$�\+Λц=�S�S����dE���j�qt�����`kY|EX'�;1���dܶw4J�Z�F�*��EnѴ��5���w�g��^�EDy�lZv��G��>��J��΂��%A+]��&LA��.&1����;Be`��5��X��TV/�ž�;6��*�R�p��w�"���r��/9�-y4-Ѓ#y`��-c�b7o5�jXm (�ࠊwı!!G�K�\6a��2;X�dF��a$K2@�y�S�]�"V�6Dw:$�)��)%��+w�}~f����s~�|�Uud�ev���L:��s�+�2�GQJ5q��fFg�������t�~�E�Y�N~u,��貳-������M��Ԙ]i8rI��1f��-Z99��`䲪�9Z�Q�R�n^p�����u�����Qh��vK|�#/*ݓ���{:��6��[g#	�7��Æ���o������Cb���S�{��w$S�	ZM