BZh91AY&SY#03� _�Px���������P9�� �@Q�BI0�OHyA�0��41�P���a2dɑ��4�# C ��A"�z�OQ�i4�h��14`LM&L�LM2100	 Ԟ	�S�#E==SA�M d��i�* �MƐ���"�S��I����3��_AV� `��PI�!4m��0x�Uad�lB�@^��>L���%Ԛ��r���xg�nx�H�:��k������w5"J�OD��8êōbQj�Q��,���i��a���[]C��@j�-+ȋ�ҟ�d�7�"Xt����&���@�������!8qԋ�������ǷȰ�!%5u�Ht�r(T�+߱�#?��fP�޼hNN�N��d�#�������Y�s��ÃȉB��!Ga�&R�%�}��wAB��%�yx%�#������iD�U��A�V���0�ƄcX�	����e��56
/��v���ʬg&��#BJ̑�2��d�,���K�٧2N^��p�FyaΓ0�N�vN�B�β�u��8��5J����+咞�u�M`�Ze��d�bB�𐄄%�$�P(�ϗ�v�0�&#��9d�
��#�#uC�$����7 ̡$zI�G'(j2�Cm*�$)qR�s ��Ą��S�g`a��d��P�������O4���k���O��-�+�x�xc�+�wf$���T�KA��3�a�f�>A�� ���Q�u�� �
Li�yn�^o!��_pt��������!����( Õ��'
��I
��H���b��҂߳I���o>4;�TL��༤\6��f�o��A�[��@�ku�Ճ;�ÿ�Cvj��P�<#&��� d�4�r0k�VЧe�vV�p3˙cR���1(��
�G�X=������R
��z����)���d�A���$������!v��[j��Jh[[^9Y���b�b	���E�	�3^{C@��Z��z5-m$x^�<�4fW������T��*�K��B����Q��`�	�D��+�
Fƈ��l���a��:�`UEI�*9PJ&Ȁ��Aͽ	엠B�zM"9�x�8?l��#"�8N��_��}��4&z��AbI	��&��3��!bB�犼���.�w��`�PXm:�fY 4�����_�Pf��t����0�gH�5P����U0��!��+Hh�e���H-a�v���Q@Ȗ�VH��ea��d�����`���ŁQ-rJ� <xhmy�-w��F�`��QY�<��H�
fp 