BZh91AY&SYG�W� �߀Px����������P~rm�N
  ���i��S�S#F�1��4�M&�        %=D�?T� ɲ� =@h  s F	�0M`�L$H �4G���6$�<�mOS@ FS�j&��� (�!(?��9�hRLbI���M��p�UC(�f)�� �d.��5�i�˽�ٍn<�޻�8��ejJ'����9Lb��a)M"��5M�E�򬌾ϐx��B�, �s�_q��a$�Y��YB#���jkk��0���9�
 |�E�}��&�+�����*6sȰ�GN����;�i�둪��ddB��6*)Ay �:{�Q���� �^E��й���kј����)��k�
�Ƌ��K�@*HP�m���bV�W"��VP*P!K�_I�XJ_*�R��!J���Fu��5�,A{5Ђ��1����Z�K�j��"� �!�	���\��'O{6��ڭa���L��!����P�(��UX��O�`�Dm��S�@�d�gW���%�>�x\Lͭ��	��JHȤ�#UvR�*B�D��PP!,k̛��
���Գ�StGb:֤���px���L�x�#��Ŗ����Y�#>#�,[	fk7�Iͻ"Naa���`5�N/�kH��$�zAP]/�̹��^iB+�z�P4&c*�f�B��hW��'�j���%�*������36��ئ��C7u��A�[ڒz��m�*��m:����s!C��h�2�F�D�K��_�+��.�r��p3��Xb�gcLcm�	�F��w�gX���w�L��2��s���O% ��P��Mz�"�dp�E�'�@6�P�K��f)!T���qx�;�W�fܰ79��nb �����k�>b�k�$����g`Jt�����q�%�s�1P`b���-,�t�G�$XG��L��ɎDAG�E(��� nsS�AI���"l��g��sB{��A�h)��L�i��u�߉�`����A���8�A�hL��v����`4;�N��h&y�,:���+OUB��i�4�d�4�2�Dǈ�|ѡA���V[�KŬ���MI��PAR��p00CP)5�u��m��$\4M�Ye%*����F���F�G͑�I�wi�o�$Xp�/*#^d�#L�>�Z�7i̫m�~��4�V%����)�=:�8