BZh91AY&SY�@) I_�Px����������`?
���   �)�ڦ�G��TH�z�i��h��M4 Rjh �2h h   ��b�LFCC �#��b�LFCC �#��b�LFCC �#	4ɠ�x�O�	� Ѥڗ�B� !$�D����?��9`��p��
Hb	��_#��n�1$\4+!�a	4rjM�����q��7uW�.�'|a��>r�0��dB���H��l�f�t�%��n��r�9J9VQe%܇Γ5�G��x�i�bF#�c=�Ӽ��R(=0�q�f9�����ٳ9��3��m���t�۝{�>�#��e� 4�������W��p�϶J��R�$�o���.1�zu�¸r��� 47��9�v�*� %7!w��uV$���Vi�Q��:V$��" B�YR栩��M3�*@�����H�w���r8�{)DXD	��H8�M5|�b��q$�\;\\T
�������e^ؖD Y���X��he�Y�ا���4��T����H���$w�S��.��R��-�EU����`Ж�ۋ�t� �A�%�� �T�܃���ȇRSR&����(xF�9�4C���9d�^��+C�0��I�""QD�K�ɍNPHPO4�A aq���&0Ca{3�$U��؟{�|�߮��@���5�6�2A�_tu���1�H<����	�=�%I���xE�j\�s9ʩ�M��Ey�n*H�PTaױ,�?�� ���� W��ҤICT��)��^X�N�K�f��Y�D6�� ?�H�c#q�0�L�`l_)�!�͇ҡ���<ܒO�\�i*f����^Y�62:s�&��� ɤd��q���JB>�tV�8��,hW3�M	��cI8�P8�{�{���Yq�PP%��_�MSԠ��P��MA�8�]5��܉h���4-�����!��.�e�X�>e�j�� evk �����Uk\w�C��!	���Y���N���6P.<�y��Is�Q�Ba�9�B�����I� ���J�	�:Zc�C�"��sf��79�N�6������� "���ս	즰��S��  i^���A�`�����r���1􆱡2���,I > b�ќÉٸ �H��Ү,t�f`�o��v��t@�s&2C3�0a�S���y�A���ha�8g���X�BjN��J 3Ȉ3y��^5�Y�X�Z�H�n�ѢJ�1�T�i�=���M�����6�~�oH�q�`X�"�@{����s�Zٿ�l6A�`а�����"�(H���