BZh91AY&SY���C 
߀Px���������P�wV�:�w!��@J(ڦ	��E=F�=OP  4�*`!$�Q�F�� @�4�&�4���@   �0L@0	�h�h`b`�!�M4M(�H�h ɧꞦe6�W8Ii"2�F�!^����П���D��0%/S�~���xHkT#0��
U#Cp��B��m�l��\O�T̲��ևy;��Nu+FA��v9 5����-m��̉#Y�M��V$Vw�s.ydo~��?H�a���PGN��fɰh�I���T�]�r��ǒ7N��ĒI�͸`I�����T�8p�D-�:&;�Kj���$�5];!}�!"[4�X�G��2`V�p�L�#�Hn1�R#
]�ZDi��s�:��A5	A�Ax�Z�AK^��pNkd�F2�y�ò����I�%*2#\f|PA"qs�
P�1Fj2�I(�eYf+�n	�
Bsh�) ����4���%��KV���)n��=#��;9�
�ɥBf�C��K�E�5����jޚ���L���3V0M'���j1��\�#�������Jg/\�q�rb9�9d�*}�������E���e�[J\XI}�kp$$!
츢D1��f5�r���m�4�$U�y�Z����ฎ*%�Q�x8<"9�}h�8�ɘ`�붗��mDf��
'	��g�d�F�L�2�r�r�33�H:��O��)�V��\�-	��W?)���߉���С?�hX�mxW�ѷ�0{�Z���?G�q9|��)�����Fp�h��N�둒S��T�i#��92?��Y���D-ycV�脌�F�ɽ�Xp�rO�s��)�9��*"��`�����i���ߞ�)��4o��K"��qpf��5����8ٷi�5jp�%���~���Yq�(�=W9/=��nq����5r�afn�"�<e�����qh)/���9��q�$�Q�bŶϏI�\3�?����=�ϬO�����e}GNF�y�{E�	���ED��M/U�^�ؒf���wd\��Wv�=ceD�8\U��FQz�sDKb�V�g}<�W/��NB|��d)���.0`�|���>������η7�;{߅|�B�S?[��4^�Cz*)�,�w�P��	�������dn0�R�B����T2�E�m�m�6jt�sܙ�3�s؏Cza�-Kֽ���ͮ�Yjt7M��KC�L�y5kԹ��'�������/�K�ԍ�*���)'ܳ���5��K�r���x����>{j�Aj4Q�)iIA
b���Pc���ܑN$*%�