BZh91AY&SY��� �߀Px���������P�:�9[`U2 �Q&Sh�"b �C    �?D�l�� 4      ��&�P��� ����& �4d40	�10� H�m�)���Q�=	� L�O)y0���	(?�r̛�hR��@�5�%��	�M d��a �ũ6Њ�GÁ�џw*�H���w[Qs@�DA���X͎��y �b�!�g�9��)�6y������[g�A�&`9�d�J�q�E�ڠԂ����Q
���fj ����
�K����  �s(���� i����dYL��)wcF��7"�I-_|��� �)FV3�چi��F�M�SR���*������[ak���e�z�5��	xn� �
�U����-�h$�D� ��<��15h�ji�w�bO,�h����
�au�I6����Zo��<�&�)��������c���CAw�l����5rZ]���xav^II����G�Z\��bF		��b����A0�-��5\�( ���,�1t3;��2�|�7s���ƟJ��Y#I���4_N�G��)�&����GY&k�̎��&D�d�0�R�WB&����H~G��.�A�� ��/:܌7��ۥ@��%�x޼�[���Q.d��3Y�@�����x�D�L�j(�AȷRI�P%Z��ꩻ�O�.��
L�P����T�A�^���0k,R��T����������"��Cm�&6�0(����^�s�H.	,*F��q�t����AQ$�Q%�I����i6�$�N�h�腩���hP�8Ƙ�I��hO�>�PV��,T̸����zmkq�j3�����'�GA^��6�N�rķ
�90��(-лJۖ��X�5�o��(�a����P{^��h#�3!Z�ɢ*�P��"3m�V(O]?�ZA�s ��0>��1��\�p�7�a�}a�9�1�CHЙ]�I�$|�g�x1�n�T� �0��X�:���Wp�f
�4ݸd�2aH�&8ʕ�#�5r�x�V��r�!��X�BjO&]�
�eI�fơ��.$���RXg�MY�T��0�{02����F�Pd`kE�k)TIm���^&�K]����0h$��=���H�
���