BZh91AY&SYi_=$ X߀Px���������P^�l�p:�J"j=#S�)�`����z��j  %h�H 44    !&�jC Sj4���@@0&&�	�&L�&	����@&��iOԟ�OI�� �h��=@J� �B���~����� ɡRbXI2���|8I�KA�f368��D����f���/c�r3�Y�3�2�����������J������3�<b<π|�4�A�,0������qQȋ��Y�ėh�N�|�B���UI�,�T5訤i�K�͛�pR���
+�k)j؍Z�Э��\*N�L���	n<ar��Yŕ�-�0�jn3��F�+#)&��W�B R�	�qё����*�
0�\��A�(L��ЙY�r��p�
���$� :d�1URd�й�*H����(��¨EE��,Ů����OKYkzӨEbB�j,FV5WFX�^Ӭ61���[m��w�N�t<4��"9P�����]�l�����ᆳ2,���n�!N�R ʨPC���a���h�mF��A�_���9�ݖ�S����SL�Bw?�h�K�Q�h�����|$�_�!��亣�c͟8�ޭV-F��-,F�����IVH~6��|�I� 2K�3�1L;����^w��Z���T��hPKڒ�FL��*704_)*Й̨;�l��_$�Ơ�)^�܊�;ZY�y�n��ѐ��v_�RL�0k�4!�"&Z]*W
U��{��_a�!�)�+�IBCI�%GN�XS���l�ݢ�,.2R �Gu�=�(����C4�a �������f������4RSB��{u*[�b��L�]�пį<�4Itۂ́��@�|ԥ:u܌�Fœ�M�.�Q� ��S�>M�uǠ1(F��`bL0`NfAHn{'(Ę��� Q�yA �,�����ahN��2���D4P>���"/ݐwnBy�Β�p	��Of �� G�������7� _�i���S��	��8�Y �Ě.:�mIdK��י\Xz%�`��[�Pm:�3��ң�䉏�����n���Ew����Ȭ�jN۸$�]$�x� �q((Yu����H���r��!b7�Q	���DT�3Z�Y���$�5����ׁ�U]��dc�,�*��ܑN$W�I 