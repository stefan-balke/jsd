BZh91AY&SY���� _�Px���������Py�68��[�@	B�h�)鉔�=5 �4� C@J	��2 ��i�@ɠ  D$OT�z���d���� �� ���a2dɑ��4�# C � A4G��jL�6��OSjH  ɚ�S)H�BD$
��H���������B�L��'�p-�!\hX�ń&��Km �)H]��M}���͹�<Y�9v%�GF��������U��茰��lOƵ6��Ө>9�tʌ�#h�H����l�#�II�v�7cn�W;��4 �u�s*��H֑�%~��OX�� /�*((�t1�.B� ���\:���[��n%�@`�sBz����)��� �5�l�"�<�R5J͹w��
#R������G�+#"�b*���ď �v-[g�f&X����f!D��l�i�����(�0�0�bE���F�61�Ͷ�CB�^��hrJ^^�iIBxG.ME%��:f��c��$�D ��!��SyPU䐐aq�ej ���`SSD��v�s��.'2�9^ѓS�a������:{�!5CG8EF3���G��i�7���1iM�Ft�=xy��ĳ@kk һp�?�C帎�<y�0�B
�r��Y����t����T���Y��@��p�/��L`��fe��� ���$���[H���s9�Øvj��.8��&P��ZJ@��XE+
U#��u�|8�2W��M��cI��Vaȸ-�~ nӇ\8L��B��;M�����	��CI+�J5Ux׼.Ϥ�uF��VtB��ib��2S=��A�y���<K����V-P�yh�g9�jĂ�"J��	;�ݰ�Clv��Bzݑb\Hi ɥ9��Xn{��9�Y!f 	6hP"B���"�^�rA����JI:���H�d@E�����҄�Į`�MU e^Ԍ	�!��~��b@`1�I���0��T��=&�bHO�Hh�0���pLS5ܯ,|�ipu��5�A�恚�2CG��c�8�G��"�GH�:�ԝ�jPL$����Ű1��
��Ak\JK(T@�k�S�4�������������3��id���Z���\�^󂥯�٩�7�O����H�
۽��