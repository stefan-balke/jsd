BZh91AY&SY��� _�Px����������P�rV` J���7�jx�D�LH�&��`�1 �&	�!��L���J��1dzM��    9�#� �&���0F&"	L�i�#"cCP2 zh�1(�|��$U ]������@8Af�)���KQ�x�,�B�˰b������aBؾ`�gR�M_Z����V�����M.�P���%J�a�n`������I���hXe�GMюrSΣq����8������<��{��Z�� �͑'&`�_o�
��0cû�=�\����J�e�I,�ՑJJ�Թ�QS����*1�2��D0�5A�3��ʷ�B��D^�IA`5� �����E�kFbU���s�n��&7�QZ�H��r�"���<���Iet������61����I(@�c�S��F\CNY0*�rG.F�K�����)G$�#jJL�0w܌P�(b&XQ#*Q$�����W�D��	+�Q;f���11��@k��/M����W��bŋ��C.���O|t�صNB� �������F���$~�~�����{��Xt�G�!���~��!P= �A�@�^�Q��|�_�%��,p��2f��P�����x�"��l*�3 ���bI�"���j�8�������EN����Pʁ�3��A�"����hScI�N�s�x����=�`8ĩ�h\-�{ �^m���ȸ�)�z���k�I��!���%�GWE�!���6Y�!P�����DR�LG�P���w�Ƞt�QQ���9�ӌ1�Z߉���M$m��Ǡ��yG��Nچs�14�s�.0,T41R�Axn��1�D9 @Iђ� u�$A^�*�P�fr��B������y2=;�����8�L��"���K%�<_�%���U������%!�� �<ۄdEVK1s��@��h
��D��d�h��H�Ѽ�̍�{���������K��E/6~R�,g�ᵰ4-�� �T7Ծl	�h�+9jR���ɗy�#W��6��]�'`�؆Isb�XZen��93��ʷ��g��B��Bφ�ٙi?�w$S�	��