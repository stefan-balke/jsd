BZh91AY&SY��� �߀Px���������`\c�q�C� �L%eOi=(�=Oj2F�M��d  �? �����h     0`��`ѐ��&��BD� ��� 4   0`��`ѐ��&��E#LFC()�Tz#�4�A���?Jk,���I ]	, >N_p��~��@XHMO��q�rX��a��j�F�I�4|;M����帷�20�&�UmV-�����P+.�jۇ� oާK'#@ہ~`A}�p�wbp�&T�hۘB�Ԅ�ӎ��~�a���� V�b�i�@Н�/�����{YX��Z��Nr@�=6THHT
�"{�3�빱��S'�g�D@TPQvz�,��L��#"��GH��%���\��5z�1������4��AŨ��3��E=�4��Q6h3wOu�M5Pd��ݔ4�,� �Tv�h��I@��5�|ވei�Ԉ bQ"jtj�9g�"��hDDp���7Xņ���u��ԋ�l3m�lC`��.W�Y5.���1G �� j��zU��*>E#v��4( �:�� �0`ES���jf�@��h�(`'	��Ac)igc�de��lwW�3A\�T�x�i/�k1��61���m����v����\{H�B�;���^��6S ��H62��0���2����6�ِ�"��,��8��ʨP�*�k��ɤ61��|���Z�˱k������l��Dlc$ ͪ��He������/����GU3$�ˌe/UcZ5��77ΠW�C��ũI�2��һ�����)��H?���a��,�) � � |���0�_1�J�Ir�*�X�rF�m=&7�6�:�$1�3$���d"]�'l�4�U̹�:؍�f���2�a�SɈ9��i���t��<Y�K�3ρQj�ޠ4��i$�y5̀T��ݣ�V^�(�����|g}�x��E�:i�
��H�h�d���8�"khZ�x�3w�z�ϸ-�4c�ay�H:,�ni-\���)�<��j��f$\O����@��&N���9A�q ��JF�����oB� �G[�A;�,HHF��%�.d΀����"4d 	2Y��xoBxO`�v��@2��jJ#�yTuE��P@lM��[E�l��	��8�DR@���CG@1����AxHD�W�G��2}TA1�䁙�2#SpDG��5n�EC1ە��K-"�ʨ��IE�ә1 ��*`���5tK�ˬi�A�F������HD��>
=�"�W��kI�� uf`��Q��Q"��7��2���oS��ݗ��M9����"�(H
wQ 