BZh91AY&SY�p�� �߀Px����������P��]Sc�M%bj�	�(Ѡ4=A��h h �S4L& �   	�DM���ɨ�CM�  ��& �4d40	�10T�M6�lM54�$Ɠ�di� �bj_$WL��A�#(��W���*�,�T �B�` d��~���!�`��!����D	DO��k��j����f�MT���|�!D�?��H�	S���-�R6�A�����J��ƍ�Ӭ:t�1��0$�+\�5"�NDRMx{��-�ƹe}�%K:�@	c�.�HW5��=�]8�1�vH�����1�bY���A�B��T���$I�Q��M5�5�R�Sc��&��
�#]w�Mf�rn�[mY�<�)C�a�K8�$�X��4�%�`@V�aiR�]%YJq%@���E�h"�
�[-A���2��%9ԇ#��Z�W�M�y�a��4��42І�����8�e!�k��{��\�����ɦؓA.ы;������7��m�4�9(���\�d;�JJ@���j(�.hw�q�Nvj�.QXCw�E�D��$�S#d0����`2�AX�! �ם��"�J��K��fe����8*8r�Cǩ�3ʗ�R�e0���`�A��a �	Bk�,�MH(��c��[�X�dJa�Ng�P1(G��qZ f�R���o��F��!����O-w��yy�yKB���-P�o�{���I�HzP�Ftm{�0��gE�ݢ_)�6�8����Y�1�I=���堸�-�Ż�xB�y���Úu5d��3Ri!��!�Y�ׅ7#�͗Ft8��`m�����m��8�,k[����]�2���s46K�R��g��~�e~�b�������yG��׏y���m�Ŗ�Վz	b���G�Ըi����h��t�X�Msm"�X����jW�qφ���3�����WK�*:�v��WX����9Y-�L5���_sa������]�ab��@�H��yC%Y"C ��{+*��_��������mM�#�|J����k�/yfmi,�.�V�כt�N�5���eM�:oWaΨ�K4x���кB���Tj)F��r����Y>���x�C�#�Y��V�*\�I�sZ�z�:m��M�u�6�t�y#7�dU��k, ��H �4��6�8�
��`qţNK��T;j��c3;޵a�1c-͌��R6|�~�꒤}k8v6�j�s&�����p�c��ET�:&e���ǅhmQP��+�.�p�!.�`