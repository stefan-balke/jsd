BZh91AY&SY�"nz x߀Px���������`_z�'�  �h�='�HdѦA����&@ 4 jz�H  L & 	� � �`�2��Jz���@��4 �  �`�1 �&	�!��L���h�d�&�z!?SSh��=51��� |` ��$+������F�@SP��D%1�>��))�4$\4+X��:ڔ�	Y=�Cn�'����e�y�Y�[���iw&�lxΒ�����|Ϊ�����C��4��;]eJh�u���}����|\�ՙ�a"�,.1�p���x��L�ctAI���q�20�X�S��0-�����4&3%����JNQ3ԙB�g�x����cm1۫���!+��p�˜��d&L��5��N�P����W1���8��`M��&�p����$��ADV2ƭ�1���5���R)�׆ab rMv�$�&̓M���i�84�K0j*�cr�=��Aw2�K�ZˠCpf��
���A+"`��E%(�[@�Y�kV�ʚ�����T�-!X9�L.C3%H��;YH����!��D$4#�1�֨IG8Zװ- �.n��ƣbk,���S��k:י�t�D^B�� �v�N�wj#�i.E]Sۢjh��^
�DEc&1CwE�\P���`�R�,(�I8$%�8RĔ3�"KΊ
%����	����a)C��Gm��[f���;;Bf���ц��C*��-�P{��pw}Ɋ � O]�=����{T��:2����g>�����	�2�$4L��Nm���g�y|�LF�_0�{���B�pB��y\�ˡ}FY�%��	�`��I/b�gځA3cZ�D�L�k(�S ���Вy��l��@�i,��8�Pkd"��/��Q$�!��4!��&_�&J�%��j��<:L���@؛m�1(rd}�@=�k%�*b��-�h|~T����,�"K�I��7=}an[I�T��4VtB����Qqu3�L���?'�}�u��d�WfY0�x��ֻ�q!�2��#Uv$�n��R�#�l2�^s�:	mIT`h&g�NF��7Lg(�LI�]*H&@�X�D�>'���EB�f�G9�&�h�zʠ�=�P�<hO^���$��T*��b~�$1R���M���:7A��=@����1���2���	 �	&��c޳�bIi	�I3�J���7��8�h�ciށ����"C��m��Fkٻ0����,��$XN�5'u��J��P@�Fe�0�fX�����Y`�]%%z/ZI� a0��]�]�#'��H;�9��AsZJE��yPd�6��}8�mxU,��f#A���]�붟���)��s�