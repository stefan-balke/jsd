BZh91AY&SY<�; ;_�Px���������P>q`B�J�$�
x�Q�z��Hi�F� ����&L�20�&�db``� �� ���#�P   4 sbh0�2d��`�i���!�H�"���ꞧ���S�@ 4�4����! TH$�?����"&iB� �B�Ц	�k��M���B�hVtL���-�3�n��SZ��tO-¯�Q#����6;Gӂ)�T�I��J��fuf������IQ90ht���
�Zo4���s�v�O�#��s�I"���J��A���S)���E�&�1����_HE�p��I-YR$P�+)�ЧZ�%_x�
��z �� �auLB�J�C4��?+m%����V])fX�"��.�k�w����E�X9͂��U�KS+�嫖ViL��B��to��N�"�I�h�;��!	K	$��Ag���I��uF��HU|$r�n�)a���V&e!G4ʹr*M�D��e!���Ē��I�� ��#�D���o�r�/S��h4���}E7p�c٤�x�����݄��}��t�ShZD�7���R�!C���hZ�h蚕R��̰1�_��!!��}��a�4��y��+�l�$0��B���F,�|�7�6� �`�f���>%��OMU���U������f���E	r���ApgZhv�5�)XRU"��6·<yVnp!�8ġװ,���h�����>g�~?�5jL.26�]đ�Tv�@�od��CEgD-��ۑE��H��(v3y��4|�����%~���ז��<kZ�r��Ұ�!������,W�|��� �ĲF�KJs5a��9F�r a&�t2	
U�����G�u�*	��=�.(X�!���T&��e�:pB{�m�;������"C�/u�# �9N�G�7�	��5���A�B|@�M���Ѽ���yjW�;�7�3
	E�l�"D",�'���/�Q����*�+�2�L�"��Rw��(
�3H�p3Q�h�P�qR��I_q ��.E%�
EP0�#u�siy���Lq���6�E��1T�� ˇ� �u-������4F&�~�����ܑN$�N�