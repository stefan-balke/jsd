BZh91AY&SY�4c (߀Px���������`?ض���  ����ѵM��ԍ4=F����F�h ��i* i    4 ���a2dɑ��4�# C �)��L�Q�     9�14L�2da0M4����$H�	�)���i�z@ ��zLƂ�A�	$*��p$@��|�!���ciM%0k�?�6�^UTE�IY�����9(�E��ѿK��N�lȅ~
��9�-ݭ��DC����SxO�K�\ZE�Ӄ"�D�$�z��+bU�P(۸X��|���y��eFX���H���83�"P�d�<2�A�jx�&����i���G�A��j�m�ݼ<����U� 4���8u �#h���\`@�|�G>�2�JB���X�3�h���� ��������ٺ�Zx�6�Q8�ʴL�r�����tB�.ĺ�}��*�
#0K��'ͦ�6�8wK�y"`*�c�a��bo�3 >2�VԢ�%0B�zh"a��G�-f�`-Q�U"�C��qĘ��2���N޴��X�0���鉑��q*%aa��0���
2�Q��>�RFAUj|�gYl=J4���ԭ֓NM|�X�0�A�	'b[m�� ��8���]�9��nĨ���ō�C�"��D�T �	)>Jb�P���@!ʬ��H�$Na��TA\�����0�A;�H$!�l�ɀ�@EP���*���yQ%��xl�@�fPxi��;[�}o�8�%c�N����(5\�@/N�4翋�H��u��Ui�Y���^m���	ԤP��-��0�B[�U�{����0@P����%;��כX���2H4I��gKg@y������*�� =�TI�9�74W�܊&!�ʇŲ<wM�DR��4�,��t�v��B(K��
$�\�b8��5�R��R=V��cȉ��/*�g`���c�%�8���[����a���*b��*|R�q�w�]�� 9�0�i��8�=�l�L�g�dB+:!m}�7\�Ц�	�A�}1������6 /ε�  #��?M��z�j�ey�ˈM-L/{b��q����,v6�XbT�Y
� F%C;sY�nz'(��I�+2�
�T�P�غc�C�"�	U��Xs���&�����l�w���Oe5���!Du��E��
C��OF���#z�2	����17��Hk4�g�,Ks "w��&��c9�w ��d�,u����&�:�A�恜x�Ɣ�"C�15���,3v볊Њ�0N�bu	�;��P �����f!�g���,,a���놗QIi�D5Z�<Iu4�?G���h<H:=d�&`��ؕ
��X0��9x@|kAU5�����ۨ�`��#U1�W���"�(H��1�