BZh91AY&SY|��> *߀Px����������Pr\��X  U6�����i�44h�� ���j��(� �4 4    	L�2T�jI��{Td22h�����& �4d40	�10� ��� ���I<��b2 �����@>H��Q ,I }�?�r4$�!Z��0L�_C�7D|�,�B�e�8�&F��6����>Y�U�ՖJ�\{҉V��CN��Ybȓ:��$��=�"�|ǯ���e��Te�r����q#Bx�Ki�����HӦ~����@
���J$
��/�4bw�)m׏�]����BP��AƠ��o.׾�Z�̎x(���61����OR�@�^�^�*;����HJ��.�8�d�*���yU��%�BE��+f@*(B��A{��$%yZ�gbZ���.
#�!�4��@���V���.XV�T���.�x���7�m��Р���szC�$qyF��HU{�9r7U�^�rD��)*RB�p�#�R �D�h1�2�I! ������$$Pb��êe;I����n˷G�4iGl�zU��N� ���,�a��m�?W�;Y�6���H�]�}\Gr�L�diG��Y��Nd�m�7o��r��|�Y�/�B�����)�`2Pń��^��о�,ޒ��
���x�K��<(706/���3"����園Na�l��Y�uc�vB�&B(q��ڠ�@9�\�&;]+
U#�Ί܇>�K�~�11(sdy@`n}a��diT���h~_iҘ0\�d�Q$_Tq]5��m&A�P�IM'ז`^�zɜ��_�.�,Վ� Y�Z�PμrG�k^[v!�B��Z����� ��_8����Zt��n��CI���V��\M!Z@9�P"A2J�r"i|G�Bv3p�9�&�h�v�����!�nBz��Z�u�@�ۂG��<����M�� t�A��v�����hL��s����@	��a���X��3����=&`����v�g��"C�B�.��e�~qV[C}�q���MI緁@U-��!��@\56��3g�H,�b�RX��"�H%����������b=�>cPf`d),�R�H�n��uͮ�j���vbq!H��[����ܑN$%�O�