BZh91AY&SYޖ� �_�Py����������`�z�ݻ�1��4�����P�F�I�@� @ M�SR4 44     2i�# `F&��4� �S�$T�S�4���h� �dɦ�L����0Fh� I @4�C)��6OT��i�&FF�����"�I�D�(%����*�؂8�&) a��ȀJc�pZ�G�&�DȦTZ�Z<*_qj-h�E�1ھ0Yr�η�]U$ح�gefV�p��,�>C�@�Mt�OGVq��4vh���wB�����QJ����j��o�;6~Go�~ӑ��#T6��ahv�$d4#�h;
��!^;P�7ֺ��$�jۦ��I���'l��:�ru��ݪr�D����,����� XE�h����t�[LRL�=
>�RS��A4Q�1��L��H���<4ԈזDٖ	�Q�'n���85�5��7��A�T$(�ZIeetX�D�����1ja@�35���D������gK �oX�l��2H](l �4�r��W.��.(��2-�˻�t���T(V$��FP�gD̼4��ʌ��,:,1��D��;UcDV0"�#�N�N&���Uh�	!�<�a\�R�\36��0�brv��tFmC;]gD�n�+k5t��KLBS(��X�%���`$H����D�o`��t�l�jJ q;�MM7W���gm�T�<L"�͕)S9��h�K��*1)�ᨈ�c��IzPPP!,u#W.@���7��?��0�#-�����x��yۦ� ࡷ�^��@��D|Fw�T�DE���<�1]91��z�6$�@�A �9��0���bTEi��$>�����xO��-��0iइ��,n<�^�^�[x��bw�'�h_ˤ�����I�LdN������`a%;(qU~�L�R���b{|�e���\��`]�:4��J��N�����RκZ-�Ѯ�u0
`9�9ʒJ]�E5[m.ķ���늲����l��R�*ٰ:p21�+��������^�0]�s��g~r�$;��p�/�*��|�&>G�̽q�[(�l��k�Ǳ��3�ϥ{�M_���.��8$4k�U��]���jVx��\"�dۅ�&�)����GF�*��^�y��݉0Pڼ�P_{3U_��غ"j,,\眲./Xq��D�,�'C(� ���l�E��ɂ]Q���E���2xr�]z[��wq0��"ʑ�+d}:[\&Ȱ��g#�#7o�
��y�fK�����QMe�m|ܒ��sK'��h;ӻF�T�P�wr劇�����F
�7$詿��)˷���ю���u:es%��˫N���\������Z����x�4��%���7F��B�וl�e����ƻ3q�)�gw�s����/d�51�u�go��uS��1ѣƛ٭�ka�w$S�	�j�