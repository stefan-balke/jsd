BZh91AY&SY�xQ� �߀py���������P�:"�c�L�I$b�Ҟ5� @ hi��4�U4` L      ��JO$�SA��z��z�  @2i�# `F&��4� �D�&�ħ�z�LS��6� 4���HL�� T$\� @����b�<�Z��&$2Mx�	�pw�h��0�4v�B�lh����9����k�u�ŭf�-+4VzA��C�a��x�ŧBD�N�s�z�8�<�_��:6�2�,H�s�9/ �O
����KA�F5�h���阄����4��%�ص��\��_��.������!a�� B�����#� �"5ωgI	�1�7��	��0�T'*�9,��H�/nH�"5d�-+5�3�97V� 4J��	�m���i���"hi1� ����MN�ST�+%����Pf��V����Dc0RS!BP�V�@ޔ'W6(.�Z����	�����L�k�3�A�M��a��d���G�ȁt�Z��ɄH�ʎW2S4�A�61����m�4��p���m�9d�
��\�փ&%F,�BcB�]b�Sz5P�n�%C��B*Xe$2����@�[���a���hs�f���r��K$�0@Ō+�I���Ek\�F���[��ƢSC�5`�Sxϖ5+걈�	��D9�zF@S����V$]�-�־���R�0����@<�Q�e+� b$Du�2E���1���KϬVI�#��k���TL�`YxY)�&C6(ݬ��}�'�U���UE�#�uj��A����3j��,��4!�DL�)XR�G�M������Yi�����E�`X+�`��F��\d�(
�=����� `Ď<f	���9���z��v�Rdʡ����lu���UoT��g a���LI
&,�u&VX��텦�<jc�y��CFА-�H���`4q+�>��e�1*Fe�*�
�
s5���;��Qp@i	7�C ����B����H丂�0�F�T`���0D����f�'��č�b����C���b^bm0D��a�����L}�hL���I��R9�5��		�L��h,tE����4i
��D��c&1�D]T�"��1A��̨ͻ��*�+xex��E�
A:�)��*_!�C5V��59Jt�\H-a�t�q��P4e5?[H����mi4.��@hh5�H��^T2DݾA���mw��-w�̍D �0hW�{4S�rE8P��xQ�