BZh91AY&SY�\ X �߀Px����������P�77w@�u44k@�@�l�zBhh�L�SOD 4�4h%�=A���C@bd4 �DD���)�jPQ�h4  @`�1 �&	�!��L�����i��M���'�6�ЍA�G��M!=�!BBE����9ilB�aZ�LHd����p/��q�Y2�!!���ID0�;��a�����7�ټ���0rl�^@�e�`�=�&�6JY�h���H��&^x��E���|������014lyd3T [,�L9�]�Z��R�z&!%MZ3R�%`��J��d�ɨUebd��u�<l�&!TPQ\��b
�8�	���!5�릑�2Vd�%�>���ĝ!+*�O�$Iee׳���R�x� �A�E�cx`�(�!.�6H�J�A	2�
�sN+V r%��M7j�0#S�T%$�-J��3J�9���@�ѫ����d�ێ$���FCh�8Tt�U
�xw�jv��H\�aA�A�r�beChɆ*q��i/8��2p�Z#fH�d��p���vy����%�I$�Q1�tl�d�M�NY1��ˑ���bQ�&6�9k$J.�M�Ђ����
�"7"%�����H j6�Z�@*��$�h�٢�u�$��Kf]y��=5[��)��a5�_z{AI��I)�V��р��!*�>\y�����p�\^�C;w����������_4�@��D5L��t��^$]�������O�W�k�g6���*!x	�9S9���3s%�%d&C6u_�g�ǻK����P��Q	��!`���.�����%����L��)XD�,鮄8����J!&� q�M���^���x<���c1@P�i��
a<::(b�Mu�G=���_�1�H�h�����H��9!L�& R��<&�$�CK�!~V�� �B��4����lD��|� 9r=_Y�F�G�������mA���i`�3 �7;���B�	�P"AC��H��G�v�,�n��J�*�&��y`M��쐞�r�M�!G `��ګ�3�zx�B 8���.�6��!#���A�F��p=&�$�� �!��c'fBF4��x,�'Y�81�uX.���u@�{��L�a�BW�F�1�v�V[�u�^n���MI络��R�7�6M!�j&��ն{Xi[��,;�d�3
ݍ#��2���h^��E�;A�"E�Se�AA{Dq��ۙ��d�kf�3��0hWi3��H�
� 