BZh91AY&SY�٪ �߀Px���������`89�� J���FF� 4 �  �0L���  �M d �A�ɓ&F�L�LS"$�S�����  � ���a2dɑ��4�# C T�14'��)�=O20�z�SJ��t�ZI	"e",�|���j�KC�t�"�R�I�_UV|�I�)L��5.���ek뿹�߳u�)J줮��©R�W�C�0V�Q#����8�`��	խ�jD'��k�)�ֶMaz�Je���Ο�-���YQ���V��c2�F�ZI)��J�j[{کV�RQ�iW����V�גLL����%JLsZ�3l�uF_���g���J)Z7|;�o�ўpӡ-w���M�^U��*]8�����o:��U�:s���/9f�&���9�I-�PgȘ�	�4bĈ�u�q�A���ɘ�6FT� ��ƍYE8�:�Xb�4b��.Q(�^�{����%���g/�-�*�YKX���dh�䢂��b'+U�E}s�������CcEA�EF�fliQ��d��Q����A�<X�6��4VK}<;�j�"(Y���M���iVj�0C0���\d�y��Q�6����\4)%�i�I$,�7�!	KRI$�P �r�{�����CNY 
Ͻ#�#uj�2�Q@�4��h:��d��P���6!(�ěi1�#�!�Ơ�V3�8�}�PBA�:r�����_q��]ޡ$�.g��$�%��TT��^q����a��-r��;ETJ��19��^��P��j�)]q!P+�>���%D�e�.��v��zgW������3mP?rб������nչ30=�.�ˇ�>؆�	�TˢI����G�X�K�ۜ��)N�8O+�Q)job|=t�ϓ/4���]�9f�1��+5�f�eeR���`��E�j`��N�Q�E�NK4�9Z]���ӷQVS�;&��Β�U[k	׼��̯x�W�Nss;�`�1]����Û�Q@�q�t�̨��<;�������NEF7_�z8qa8���0j`�)��?9��Ϳ�[�3��-�}w��q������������~�y����4;M-��Ή&J�5���1�U��}��|DA�0I�d2	
�wCccP�rZ �bH�����P\<E��Q\v���D��ہ��x��V��ԏ�߆cݭ��Xvz���>��ޫ��s*%0��qt�Ve�4=��Ш�)G/?@3�f�������zn��6&
�ZaN�*R�*<�QR�j�V�F��rb�GW-i��-69es%��˫>�� Ţ�K��J������e�2�,�l.�f�it�m��_Ƥl�W�z���,��}���s3�ic5�gOU��V����e������EDѭ�χ�rE8P��٪