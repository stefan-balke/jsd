BZh91AY&SYNT;\ �_�Py���������P�껳gSU�d:$�M��OM51#F&�4 4dh4�1M4T�1P�h���&�C@$B%=OA'���L��M  ��dɦ�L����0Fh� 	SH���h�MQ➦�4��1 ���f(@�RH�!Y0K[H% q��=�Q�$~�F%#R%���u���%�1*��D h����V_���tu�ڝ�"�ܖI�����X���Wh��#nvO�\C�X}+�1��������ċ�N�ɜ�$�!�D�J8��1;Q�}/*�Hе<�"jH%ȸ�Xd�rB�"�(�3�9ᢜ�G�D&L��w���D�	5�%<T�!g��EEYJ�s�|�[�c}�Ὁ�L�KI6�����9UHʨ�4�8�n����>��G���\�@ �*��C9J��1L$�,f&��ͭ�+�F�`M.r�aGl�P�(ZZ����2�M^,�t�T]�4xڹ�8��c:��k4ZP�(D�zO�wG�썌lczX�m��A'n�9��ɥ%$;�%蒢��׹w�jHe�S���V��
m,���.Rd4cdV2HH0��y3q��m�&k���}n��!N����9����n��x��HËCc�kj��5y[ }BP��%,�ZsFD57 >�p؆lڃ�s��R�ߴޓh4A	���)�%�F;�j����wr0�ѐ�d�BR�r�8��2%�U/�%�#�ѕ�ǴuN����65��
$̘�W�TM���3l�<�����=�o|.li9i�:W!V���E	p�0�CTA�:@3�"���&ׅTG����!�k���αg��^P�5�B����\��� ԭ4�
�XNde���t��[��%x���io�*$�FGya#�h���`�'۷Ű4��p�����r�T�B������d�3!��V��5g��v�*���ͨ\;���>���]9�/��-�&"�h�t�AXnzg(���fa�&�QBD�;�M�� ��E�\6Q7gXf�.%-9�J)�:�j<�	>m�!q7 ��\x\!��mC�ir�r�e�z���1&Sy�bR���.Hhކ4tvs!T&�3ļ-*f:΢�t�+`Lm3:m2!�N�E��$g�M&ݽ7�C�8 \cY'`MI۟"�VtrМ�5+α�!x� Ĩs��h��V�H�RZ��l[%�	��Wy<�0i4/AWZ-b6$H��g,|��t�F��6�W7���#Z`ĭ�`���H�
	ʇk�