BZh91AY&SYQ��� �߀Px����������P�s�`R㎻��A(��j{ML4i��ODh4  ����z���     Jz�F����L��6FSA�b=#�i�� � �`�2��*I ��C(�M0OQ� 4M5/�+���A�#(��W����渟�D���
]S�w�U��x4*%���00jb�	� �d,�<F�m��:4�WyĖ�:R�X'��On�f �ݜqgj�2�$�/���ݹ��.W<�#�l�b0A�R�]4�ޱ�v�]�ζ_冹��V��L�䉁��g2�1>J{�����1�s�Ӕ�B�a0���kC��H��xk\�S$�i1ܵJ�jwR) �o�l^-���a�����<p�x�,YEm���<H�b�G�U��$�1j*�(�M��v�Tr,|8,-S�i�%�k�jz&��Y1����Y��[(��n>\�}S�5�h9y�;m��i��b�%�5��΋W�#m���h�qđ)�����7D\U��	$�˨3Q���K��ܑ/%�Z�,B�T���b�+�gI4����Hq�NJf:��4�!j�K��PP!,gșP X,���ut3��x�ѿ[~��������:|��m��Cn
T
h����BW�|xm�R�Ĺ2�*�"�F.&C�/��Ǚ�Eh��&�	R���̌�����(X�j|����	��Rа�O��_��{���$�Դ��zP����w�	)�C��e/��Z�|1>�Es�g{3.-]��$,�A��L�%�`��w*�B�'*r�$R�(���u�T]y<��� dO͋��Y=,0��C;F#=!7 ��<�.+
		�! ���qO4�Huu`�Jia<k���������E�1DT&RPJ�-��% ��D�"0���}`��:g��@�#��`+q&��QgkZ�lAD�����C���
��x���c%�d�Cb�]"�یmU~��Z�V.xw��@H�H�wzǦb�@���vUa|�&	uFG{"-}-b�����tD���C��/�ؒʑ���dy6�OŲ.>���'����z���Sǡ��t�u���R��������42f�]�Rhvdi��U+S��<�mִ^��oE��S?����-'Q��;��ľ]Zur`�-7,��S���ԩd���'Y���	��*�ۡ��7�����L������p�*GԳ������E���SS$n�,��c��T�:fe���ʆ�N����)��/�