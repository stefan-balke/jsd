BZh91AY&SY^�x� �_�Py����������P��;��s�F� ��i�?)�H�@�     i�#QH��M  �  HJb4���4��j~�f�4hi�hy!�8ɓM0�14`� Ѧ 
���BM�&I�)�=C 44d�%��D��KИ�,B����V�"�b���D�,�)��:�@����0�h�j�HČH=�Mܻ{۲���S���6�mv�kt�������Bo�)�����}�`Ix}�0�Wd�UC(e"����s�N��S�� ��BQ%�"ǩ&6X��pI�2�u�����z�V{��e���&'wR��Qp�d��X�����G��zBi����<�8�l\Av��K^q�����]t����3��dLAP	�C���-��a،���̢#@u0�&k+J�Gu�F�cl�C$(4�Hig� Ep��2\g�C�4���q��,��
IW7v�D��n�0+�.X+� ��D��I`L��p��.p(F�qK/&*�F��(Ц�d��QqRs�۬�#\�:��*1񱗽FS�<�X����:NQ���okm���(C�ŹýB��ʅ v�J�I��W#�㪃i��E���"�`�Fӏ�Q�YI�CQ��2Ε��c��md�M��s͝�L�_��ƿ 4;�|='����>�n]U�e�χ�' ��n��@��_�zo0ʰEж|̇0Ցb�ݶ�n$����3��|,�Df�*D�B�Y��]�Nܹ��`o)l,��e�x'�M�2K��Y�ҟ�M�}�a,��#l�fH�1��g����u��RO��W�zb�8���[�P�Y,s�\�Y,��LV��n��e�]OC9����8V�(6��REY�|��ba֯@�WF}�33d�,/[�򝾻�]�¥�H�V��J.�%����l;������EFW_uvn޾o5˧�s�HJ����*�Z�
|UZ
�M���D��X��I�l�У�m�"yz�H��_�V���m�wA����R.��^7�ܟB��@�w�(.X�����d��Wgp�yd��aSEù�IeԢ�����'oLJ�ͶD�rK�65��Y#�݄��<����-�{æs8�-W�ܨ���yLV�hY߉�i,Q���"b]��;��3S�r��Ѩ�U*�S�-R��g6������nt�Sv�u�Fϋ���q�k2�K��i˓	V�����f��%K�L���1՚i�:�UU���k&0�5y�J��ʸko�*Fǝk��z��ZŶh`�vŎ���j���/�޺lT9�TM3��H�
��@