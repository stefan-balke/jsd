BZh91AY&SYXe� h߀Px���������P^r(�Y 	B�~�5G��~�h�C�P���@C@`LM&L�LM2100	L�����di��CF���h@9�14L�2da0M4����$HI��OH���  cM'�Ě� $��H,��@�]ߨ�d%�hRJ`�_0>m��$��Y!A�c�IA�V�)�6�|�z��,�;؅dܔH�<kFu�^1X�dEkT�*z�p��h�V_6��˷ȩ�/5��,H2M2f$I56㓜�"1Z��HBxa|�U����3K�����@0c�o�=�NcP��ۨ�F��(�J�DŜv^��Z��Wؾ(��F��:זB�u��e�eX���� �)�m7bm�ԩ�й]1���SC�
�Z���)�&L��2�:jp�����⬾Ғs�EyX���X��uW*�����Q���s�wS!��I��q���m��==��ᘎ=NFH
��#�#rYF��$���L]�je1�%m&�C��̊R���y$$5MU�DH��=t3�U���&w)5�h���(x�yg��q�	��i�:;�&4L�Ӏ?a�h��/)�Ae8n�դi����*S2��ؔd(GпI�0~7X\�>@3� 0j���A�P�
2r�qg%�2�^��н�ћO��f��C!�
���dw�$�t	V��UZn����vj��P�,#�T�	��0k�VЧb=�ꭐ�g"�j�@!��B�F��W�~�5�~��\h�(	�'�=�����D��t�6^bH�Tu�+��s� �T4RSB��7[�53�����}�/av�y�@:0�mh  #%�1�9��]P�JUH: ֗ �m��.��B���4�X��05�	���������$͖�V�������X1	�6�`*��@���6����B{)��8�`33ך�#�^�`��n2��ո� 3;$?(k)�u�Đ�����=��4	�3�Eyc��Pr�dNhǈ�f�Ib�-���ͻ�f*�+�e�38ZE�'P�7~J T�C �s,�!�A��v�j_���YIj�D4x)�4��^���&#������ �cb��6�D����1mw�-w��$ �0hXfy��.�p� ��j: