BZh91AY&SY��� �_�Px���������P��F2�� S!@%����L��jF�d���&@�&�jzF�@h�     	�2HFF@ �   9�14L�2da0M4����$HCA4'�6���@�M2dzM��'�I
 �$f� ���{�[��A��2hTbC)�������`e�@�9�)CI��-�OFt��$
��iU1DC�'U!B{fx�p�J��x�vPAll��2�1�e`�q��84@��m�*2ČG:Fk�3'��L�B�KdۉeL^y�����@����$*��|�/zcYP8n�T+���Ġv	0c�_��x��4Z�.}qJ\��a2��K�b�q���+�(��»�겑%�p^F����h陶<���C.��3�Rm��զa�D���:���,�F"Tj�
E	A�\�@hH�`�X�)��TL_2�5�����;�U����Zm��jkU��(�H˖&�<���*�jR���ׁI��I����$��)Fر�q�|F����7�m��H�;����%��G�V��)��ʹf
t򹂥��C91t�1J���wJ�Ȝ! �a�2���
�"�;Դ�
*�R�>���FP�؆׍��#:� �=t���?�hqH����Җ�,J�Y��~�W2�f���D[Y9�s�����c�2d$��7��޻� ��A�i���A�h;���2Ӑ d.� �k���Ey/��qIyy� �{�"f�7킢e�/����f�z��4��b�;Zw`U��s���g,��.Y��T����0C:DL��)T�uW:�r,iW����m�I�%;�^�� ���d�����Ab�|�X~>��`Ď��K��:*�]u���ɐeTnEgD-��V(�%R��lw�V�6��$D�!;�I�`0#B��3�Uk^���ѥ`��7�=������l6P3`���� ,01&4��`e�e�善H
:��PY����{	��0��ј�Y�DI���Xd@Fsv"��B{)�H�:0��iIj&@����ہq� ޯ	L��O!�z��>��4&W��8��$��":��|�����L��^X�;���8�y��,06��f����%"�0j�n�t�o�"�Æag8ZE��&���Ġ�S4��ֳB���o*.�y ��#���D聆/B�SH��{��ZL�_���6�cd٘�F2Do���{k�7�Z�ᚋ�A�m �9�O�]��BC�$