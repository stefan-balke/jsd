BZh91AY&SY�AZf �߀Pxg���������P����C�1d ��zޡ��m#FC�4��@��h� 522bTl�       ��?Q��Q�@=F�  �42d�b`ɂd ф``
�@�ƨ�i�b������ �S�q-!?HQ �!#B��B����Ėr@�1�AbC)���������a4|-U� � n��×�����=��V_S݁�Aљ�x�<����#j*7H�S�ĺv�T��2��R*��]������&Q.�k"���x;�����tǦj��9����I�&Z0�H�(�EP��qf"��� M��Z�� �3	�!Q݁���7^�7tߞ���Q�&�.�W�t��'U=E��ٮ\�.a�v���l���=�p�2&�p��ũhn&2[q�J��ɪ�++��7&S76�ك�r����B�Lh�}g�)���U rW`N��*�ȫ5�[�r�QJL�٪V� �T=T$�@8�7G4"j�a:Y%
�^���TZVho@@��;��.�;`��m9�1�61���m��H�=�!��C���x��B�'�D�D��C�TPک�62���V���q�dƋ�Z�c`�+V20�!{QA@�ɷ�P��32CGJ��ŕ�&�4�����g�2���O0�q�G�n���}�cL��!M�ƌ�4Ȝ�ʘ�.>$��D!V�z��fk�`���e��i#�::����?�}�i4y���-NG��n��{����R�gp���9{'z�.s�<;a�'Б�<��w�`��0t�DH��Fz���d!���O���mЖX�i<'��!��<,��2\�Ma!� �gZh{",�1��$���g��u2l�}E�HU�`��dc�W�6�ͧy�hg/K.�;����<���q�t�|c���ѻ��`��(�h��0���.^f&�{ڽ�SW��7_{F�&�*F�suŋrOƢ��,��ץ�Ŗ����K�1˄�b�%B�H߁��g���21Pڼ�D�����W�}N�Ѓ��@����(,��e���>��FC�]���0�0h�F��D����g_4Jݥ�ʑ���;v�G�����V����{��,f�^��r�S���2]$j[g@�Tt��g��FE�/xg4�t�����k/UJ�
s�r��U��[Q98[�7r�֘�1�q��9\�~%��ӫ��F-W*ʵ�V���T�808�ѧB�,�#���Ͳ�0�����z*F���RTN�]mƚ�\ɾjbL��g7�<�S�����6kCr���cӧ�]��BCii�