BZh91AY&SY��H� {߀Px����������`��l9�@�T�6)�G�=@4��z�   s F	�0M`�L5=OSDeM6�@4� d �S�(zC�#C�� ����b�LFCC �#	BL����mM�D�2 �m'�������!	QUBD������,hR�L@2M��6��`
�TVG�%D U��O��~N�J?
�x��M��c�����}ݾA��"������]Y��д��IH,����b/�b�#nbR�"`��4>A��dN4B �
����J+r�r�gH�3���T�c]�ֹ��PPc6i�@��P_�H*�m��*+;�>vh���U�@1���g���a�r̬����d�ֱ-һM �����j��1�H�n�U��q)q!�c̽A�s{�6! ��e�� �#A���8" H��ca�:�UX�T:�Sli\���2_'�&����ʴ�8t1��ĸq�_�ƥ-�3N����k�p������	|E�olEz��.���"��%�6�C7�IZ�<���P����%��c|Ξw�9WM#ew�ZW��ƙ��5
f�f��"FWE��E��h ]@����Ft��&�0�*�R,�s��p���lcx6�m  ��ggxv¼��N2,?z87xX�����5LRz.�"�'�Lcf$��RH=0e��s����a���@����]l� H(J��G2E���>�	rԱ (������i,ꞓ��ǱA�� y Iz����DN�ykSd1�b��������@�}��b@w�1ϗ���|�
�#�B1ט���ףP�A�� ��,৯�x�ٽ%��p���l<hI���ҩLd3Q��;�l�޴�+,��lhc���I��Pjd"(t_,��&P�Y&d�D0j��ҲS��g7�n�9��-1W�������mq��,1��z�� =����*b��.'�=�1�*�~z�ɫ΢h�=�{�k�3�hZ��J.@Ц���02�-�7I]8�5�gZ��|��3��,�n�1hXRHӴ@wzN 4r����U��s��PEAa�QWgPe�{8\ˠ*�wuS(�c5b�cTW�8b��nh����N�E��*"l��m�V�'��Dq��@��H��^wZ��c1D����H�d�7��広�����Ø*I 8�h��9�h��&
g�qS��u�i���8X6�3,�.��"cБ��Ƞ�{r�+!\^U�R�Qo�i����I���sB�TU��eam�$��pn��0&�T(�z����ۉ��Ľ��asA���&���� ߲�}��r�ko��F�P��_�G�w$S�	
lď0