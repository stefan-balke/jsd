BZh91AY&SY3Е� _�Px����������P歶8�0h 	D!����6�z�CF�z�� i�F���@h  � �C  BBOT��� z 4   40`��`ѐ��&��D�	�H�)�S�i�#S&� 4�f��hI�(I�IH?�����$A��Hi�P!M~���p_�	F��3F&���H�i(����0mƧDr�p,�Xb\w�c��2F�њ�y���S��+l�.���H��V%�w��&�L��K�Ŧ��� �QI��]i�@aB,FN�E!�&�qWG�A�mz��I$��UԢ�C'ԄJ%�C��Pd����}r�a�~Y�xTPQg�J�
�J,	u���Di2����|oP�Ծ	U��XA�(�����84�{a�I��s.d�����ZҤ�4ȮCd�WA�����1�S�d�$�Yŀr�B��$� %&�3م�h#�2��UEh@l"��T�Zj�j)0��b�$(.�WFe����h�H��Z�����^��w1�,m�%j�ܥbx"�e<W�Q�1�i�t�mCǧ�h61����m�8�s�C�B�p�ʅw�TJ�Ik�9u�PMCW�TqUSc@�MA��U���;,�ժi([4#[V����k�X5W����]��n���ǫ��6�)�VH4�z%����sw]k}����"�F�	Q�Iv|�sp�i���W9UB���Ȩ�*&U&�sEJK�	�LUf]�����!]�`/�!��LN��wo׸T �^u� S���:��f�)/��&TA�I��yJ��Hс��^�4C3>�ﵐA�.�$�J���Rj����5j̄E�%Ūe4M��\�0kr_Vz��hpgc�hlYڔ�,���,����߸6�)��.����e<�r�A� �!�����dtx���<��0�c:!f�3����r�U{Jf=�f����؛�Z_�͂�r ~%��1�ֻ7�-�()$�spz��0�t�����y�K�
d��9�a������@�o-A+w�âB4/q!t��B�gCpn�V�qSF�h!D��~IzN�Ouy�]'�6��Hi��U����kD������K!A�ӲC�8Йo�BĐ' 2р1�'f`,�`�}rX<���9
�B�B�i�4�d�0&6�ؖQ�����4(3=�b*�+xi�[-"��Rw�Ġ
� ���5@�׀�iP��X`���܅��H&�oN���i{�c{I�z�4�7�� R,pXB�H��4�A�݋k�pT����i��`а�]���"�(H�J� 