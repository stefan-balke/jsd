BZh91AY&SYQG�J e_�Px���������`?x  2�@��a�z�i=O(�� �  ����&L�20�&�db``9�14L�2da0M4����$$I5=
mOSOSڠ�S@ ��9�14L�2da0M4����$�e<B������  &�SD_ �RI-�DL�B����W4����
�ċ	&S_��f�6�"fXDf��$� i��9{^.�6w?k�s{���9���{n�
e���s���I+re�1�O���<'�4�M3��C���7�ؿd.2�f�P��p܆��N�eeI/G�<�8/���H�׺BY��T�����z�oy'�T���?{��%Ø�i�_G��=Kax�U���<b��Il
w��^Kvn�]>��y��k/N���n��i�{�|<�g�"�=�Ɔ��F� ��&�C��a�1�R�Y��%ԙ�0��c9��٧�XDίj�R����K�/l�EU����lm��n+�(,hՕ����m�ۖ�8g�C'	�iq�Y��)�*�E�$���-�lJ�fk����L���CB���SD��1��e��[akt�4k^�61���m��IBt�yC᤼;��B�N�ߢT�Ke���B�p�h ��j��U�2BX�(ce���ԑ�(G��b�j�Bڠ��a�p},Cbm$D�Q&#��;p��A�M��B�p�ǭ�*fP�l%ſ9�`d� @�
C�(�}�{��Ƞ�}�"Z����Y�U�{=�ԓQAm�Ab$��2���;�����w�n�$��hX�hzk�ϣ�/<
Z����$��O�L�ȹG�|1$�O�M�	N7�~R�H�����|�=&|�'��X�v�#`�i.����3:�r����]$ˤ�Z<���{",o/��`'�����z�̜V��1&�I9ɁӸ�ǵ^������f�zX�ws�~��6J)$�ܺzGF1�׏��w���EF7�}|��0�r��{��7�����6���d��kF���ŋj�;�*��{�sEF���F�x�����*:���Tn��v5�]�F*ך�/����W��k_4.;�TAb��$$# �	t�������L��K��;Z�ZŬ��7���'���5<4r��w���}^������ٍ�I���WQ�Q)�[��2]$�+urJ���R��	&�	%��;'��v3��:�M&
���B��)#"��vN�:�}�E��n���v�/ľ]Y��$���R�mi�M
��Ln��A��%̽\�J�� �9R��wT�~U�[�RTJο���C|��M�ә�l�,��ǻ�j��q�e����Cr��g��A���"�(H(�� 