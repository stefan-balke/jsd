BZh91AY&SY�W�P >߀Px����������P>꛹!������I E�*~J~����L�z�Dz ��PL�~��        ���4��4<I�CF�M  � q�&LF& L�&@F �"SF��ԓ�	��C   ��&RIؒD J� ����E�;!��%A&K_��F��@K�]�a ���U�@"qs��n��P�ر���pW@h�ZY$s�|궳m�<�G,mɜ��;+�?X���-�`ɕ�U�K�2'�yLJ�S$��f[��|��N�\�V��bE�$Bm<�Ɨ�M��L�j(�vP����d���u4Tl�唕��-
-=�q9C'Ĺֆ�,���A]�b��<m)ORwi��1���e�����sc&*q�M5{+V���A})T�(E�ԐsQ���,�@�4��З
ب-FKH�U�ǣ%�aZe��Rx�Mcc�M��CIA%��l�r�Hv&�J$���4�%�gT�!��M�X�Ò)ID����&�H�2�U&	)��H0���gI�d&`�ǣ�����v���'��e�B�C�v��9���b�۩�4��'='�*=����_TT�Fͮ^2��s5f�΁oo�M�
����6��oW�gj -���!)�����
��&TI�ֿ�����.I^�#8��*b�dB)1����	ld3A�`t�2?e�I'J«[F3���qnin�A��DT��u�T�S[��N��+���^9��|��gGr��q�m��!��^�0��} Pz�S��*Q�C�Ó�5B��a,�"Z�\ѻ22�J���A���/����c���)PZ	�̽����r�-�^�`@8�v�F�R�/}�0�X��^1-7�@2>$w��g�4VB��Z�`�� ������ܩ'y(KM��!B[�rD��T��6gT�Ҋ�*)h�xK�E���mHO4	x� C0(Gw?D��Cz �=F�_*�g6�X�C@Й=��%$���&�A��Ǽ%�U*����Z�-8,�ӭ6lP�#����%MQ��fvf��.����L���^�*%c3x��4�@���P�m\��Ɨu�KT���Tg�S��3�=9�ZMI���\�b�D�d̅�R�A�^�[]F�\�o͙ƃ@��d���.�p�!��<�