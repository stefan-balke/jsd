BZh91AY&SY� z߀Px����������`?�ݑ�ʀ  %&(�H�A��z�1P i��L�����     s F	�0M`�L4�QP	��i�CM�4�d��0`��`ѐ��&��D�	�S�MSe=M�2`  A2j& @@	*J�H�������#�*Ф4�i �5��m�	��IU��;������׬�_	t���������+��u��Y�f���#R��;�	ļF���M!MD�&�R;�f�e�R��������ʌ�q��j�Ark,4 ��)$����A��z�ɡ)��D	X6�";a0�>D�N��ն��ȕ" ����[*��V�m�a9��Y#�\(�*]�f.)"t��5I�
[�m_9П�.b1��
 w�R�P���A;�,o�(d�#�ʌ�1�g.��B��Vp��P`��Pj-�%��dG1T���d�a���#&�bM�*��0$��|�8���8� �,��I�@E�k��u��LB�4�N��9W,�(���E5��͚"�L�ːC�D�	�i��lIE�xa��e��!�ɠ�$J�7�S��he�X.Fٱ1S������,�2X�3_�mYLn����4� �%I4�헋i/,U����Q*.�bq�ݭw"e &ۤ!2�3&��T�Y4)AX9)� D�bȜ!v2�S���)��5ҵm�!EDEQ�^�_��,}�l�ً0DN��g��GGPу����0���	�r��|��iJ�:]y˚%)Ȇ5��u����/�Imbf�A�&
^��	����$�
���(	�i�{wc�U��H$�}0=:��f�^1y��Fl���(�:��J�L�m9������<��O:�[��*��t�vm5j̄E�%��epM!2]"5�R��X��Uԇ>E�����3)Ӵ,���|��b�51@P�i�'�L��H! 9r�F3QE�MnGW��Pݼ����e4,_n�r��2S^�gfL���m��mH�-�
�>H���k\�܆,VT�͢@z<gpJu���m�dX#�"�"a�B��°����H@�� 3&q���P*@�|�" ���D���Y�Ai�Ju()4T<Ő�&�.��-��B{�� :�(&,b���?������#r�/,����>��;�C�X� } k��'n��}eq*|�-E�Yqx\+�U�
�i�8p!�K��q����$5���Lf��U�V��gIX�BjN�8�H
�H��Bؘ�����T8V�,H-a��n��)�	����J}�#?���ѤĽ$���{A�)4�0*��H�~���6��KZ�ݙ�уB���]��BC��