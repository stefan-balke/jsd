BZh91AY&SYL�A� _�Px����������P��h� ��dhI!&LOTǪhh2�@�A�14Ԧ�&�     !$�oT͢O)��� @ښh`�1 �&	�!��L�����S�S�?U?Qꍩ�==&�C�h�zM6�B䒸�K"E�2������J� ���)AH%��[~�<i$�%v��Զ�,Do�c��n���vm������v2��3�Id���[[���G;�,m�oܣ�}D�ۦT�>�I��7è?�t��#�u�k�I�k�&�ʶ-����U9;�l��  ���k KGA��64���`�:|���$�
Ɂ��=N�����jȸO(�,�lDT���)^Ҫ��嬩W#�E�{�/B��6�-�;�e<U\�6�l��aH`];�X�)P�h���[[\eQ��J���YU�xP/bP\���3�!�A�֓���ե�Fhȹ<�*"\̄���9#�
md)W2�,!B��Db��j�+0"�u�3J�Y�;- B��ȵjKg���E��N�f��Vh��\Z`�Z�f�2p\��t��lc|Ͷ�C����E˸��v�	"bH�Xj㋐C���U�dK�	�xڕ�8Cf#���$�B�2F��v^I	�Q����F��5��ߪ=9_��6�z�(@3t��>�P��8��ԍ���"�ꊂ�aU�7ό�Mv�,m���C�A=�_��`[&J�[7�{r'q��Ǫuzυ�g8��uBE�cq���[�ݿV��R�s�Y.���%�y���S�M�C�	������_%1��{��r�E-M�x`v�ie���䕮�7�y�Wi<�.�ѧ@���!c�I�Ձ2�8�qLHd��`֙�|B��3�|!��'����i�i��li�r�_�0+�+�l+���.K�za����v�b�6vf$�[�ѯ:XpX�	j�Jd2*|�إx�^J��|�E�Y��iV]@��\d'X�S�q�[0�\7�&���$6���nu9��+�t�K�3��V�%�j%Q�/���4 ^Q�q�P"B���CB�ȲE�@�M�S7T�剒��e�-.���u����Bz2/���#����v�p��×e�'_tU��W[�edD�CY*3�����&��\��<L��K1�<������g�8�S"���e��TMxۊ�7�8�L-f:��Ę*�J^zq,�\�H �8n7�P*k�\:ng�	``���sIt�Sbd��k�4�&�8��],�@�NIga^I,�u��tUN��_�.om6*�TL����"�(H&a ��