BZh91AY&SY�H�\ ߀Px����������`�}�0F��=�@�S&�S@4 ����  �z ��@ �  �  s F	�0M`�L%=B�M�h4i� 4   �)5=Mhh   ���	ѠMFOHb��&A� �4�p�A�
�$-"#\(3�|��3%W�H[�f����蟼D�+�W�
ɖa �I�DU��?!ˑ��t����U�3�o����0�^5�Øol\��vgID���,���q3�"cST+7���g�mAN�[�\Ny8�f"����!���6�fPeJu�. �=E4L�Ցi���6�]i� Զ=/	�!-t�	*����ѭf��c�-s����Y��-Hi�=;��ev:"�m��V��i�ȴ�qB��(�Iͯ}nNJ]�XK�.�P
�W3N�¸�J���Qw�FZMg��욂
C��r!BD�iy�%�(F�.�J`��d֓Bg�r`�S��MA8�T�/<lqRن�!.%�	��,uzB�H]�5�
�*��0�f`gj�aMHu�Y.RFJ�,�LB��Q��t�b�$�-�|I+��Z�;:��R�,�{
���g!�݉�QZq��R�:Ћŀ���M�hF�½�QkJ��vZ!)�,��7u�n�q��B��d�["�ju�-hD��wW��r\1!���v�`u�d˓�p
"��UU���ݧ.a�H^�9��"i'X��e�U�I3Wce$��Mw"�]�K���ͦM�L��H��"���LJ1,Nl�KP� �/J�
%��aHR 5���R�y�ū>3V{u��g�@(��x�,0�"bfTSaP�O2��˄�"�c���YQ����ӿ��;�j����PCO��y���Ch�N���I#�r�ܻ���hw�]�đ�A� �4W��WD�0��L
�K�����S}[7���*X�`�|h7�6���&�d32���d|y�Na�wd��Cj�Ifsװv��B(vcN-Q$� ZI�L��4�t�/;Efyd�չ"~�5���J��"�dQr�,��5�~��d)�����q�����i�G�A���G*��ez۸����!����᷉E�5)��90����Kl�A��.�l`�|��k^���ѡii	l��$}]ǀ*����K:Xfj.%�J�Q0��'3XV�S�h&��*����AAd�X��d��L�D�uf���&�h�t* �la� w�ы�y���� ��~�K����Ö���8� ��ӂ���!��Be:�Ө)&�F�	�@A���*]J�(qְ.<�ix\.����x c��*8D��A���Pf{��a�8�I��,N�5'~E�S	C�q�B��C@Ԑp&yK+,1��_x�\�K((� 6"�i%�i|ޓsI�=d�C`\��%"�j�d�8q���ŵ�7�Z���B��B��;w�w$S�	ďU�