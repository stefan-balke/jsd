BZh91AY&SYLa�6 �߀Px����������`�y�]Ɛ@�p�і���(���O4)�(�4hѡ��F�hh�i�0R$�&e0��# C4��0L@0	�h�h`ba!#%	�i=��#ji�Q�F�d`�1 �&	�!��L����*��b�y�hh ��J��� KI!0�#)�����G	�Z	�������m�m� �4-�!4v5T��"3 Y�{������k�G!�s('�e��Äf(Ø��lٳf�"�F8_6�؆��������Y�  �Knv�;Ö^��8C9aR� 8�9<j�t��Y齒�3mU�m�J�R�-��ژ�t�pك<��7V�����Nw_�< ��
� ��:[���*�����ު�֪�Dy.=?.��F8�� *((���o�R���y�Z���]�ZY�%�eԍ��*˪�$�r�a[��m�Qv;cjA�Z��pf�ܮVVy.(�q(���-%:�+��`��	�Ia�:Cit)5n"AhX�b�TG��̦pɴ)G�f���S.RM��5�b7�f�e�FZxQ;�4�!b`ܤ�m"*�
ʶ��;b,m����ͲmM.���Ǉz��tԲ �},��
[�!a`֨j]E�x2AauF cf�� ��Q�ݑ���D�r ֐�%'D�(H��Uc��-�!�
`]�d��D�0u�r������8)0��uř�U
���2�K���#s@ROF�aYUZҬ�F�osSB�!�Uc�k��̊�"�A9��{�vUr1�7�vG�0:��HZ�[PwL����bm��T�k�Dfb�Jԓ������m��C@!㳽�h\��B���T�K��)�c`� F6����B�1�ё�"ѥZS$AM6����]\u#e �;�^`j���zR((F���C��&ѳ�M����=��tSG���Ѐ4v�y���VA��;�z&z�Ϭ��m��:=�I#];�~�x蒈�䳒I@�e ��$�I$��:�ϴ��� 9�t��b������oY灟Ƞ?�б���C�۫�08�,?�����Oj�OLQ'��5������e%9�o�9/�"������R�3{�$����F�e���=� �<<�7�P�"`�u�-` fCB�I2��0kY��YE�z��LU��{Y5���%�R
����dcޯ��9�p9�n���K��I�~�n�t�@uu`�J_;l���(�ߗ�p�\�o�
����yi��.��o����I5�P?Q�E �T�P,U��oW�ƕn�vsq�MS^�N`=]�8��a�Wu]c�7�`��w1&*ך����ڪ���k�H5D]�PY�,tHF�?a#�+,�4��ڼ�4d<�� �J+O���J�Ð�B%�ڢ׊؃,�(�ؚoK0�V	�nG��D�]oI��
��Q����@�^7;�Mݯ+A֙�bg���x@�<FPƒ�s��<'m	w:g%8��1�c��hD��es%��˫=, dֆB3�p8�PT�I��nߡA��mV�텍���/0m�T���m�W�% ����o3�p̜/��05Tѡ��*�����v�'1ࠨ$o�rE8P�La�6