BZh91AY&SY�_�� �߀Px���������P�Y�Ѹ�2r �S#T�2i�	��2d �Ѡ 	MH�M��I�d�@    �D��<�ɧ��4�z&i� �A�	���dɓ#	�i�F& �"D�d2M��h��iM2x�� =O!?Jg&��I �P ~~���h� �B�12M|E�6�sZ4*��hhbDȕ@$U�d����ʿ$�����B����r.��R�9}S
(�
W۹��,X�qWIP��;�d	���M�O<Ł^}���7Y���l��E����QigQ��;��4�-~��_+���M����誏͡��N�u�KYT�r�b��V�y��(�(�⁨���X�,���
z�5R��mR���"aZ�W)�IPD(%~���H�O%�Q`��KI�HBB�$�P(�3�x��,�i�rɅg�#�#x�Ra��6�m�#��06�0IJ�<�b-,/,�̄��5�g� ƛY���o����f��q�&os��s��K����4Ri[R��G��&�%�Q�����е��eM51���Q:����6��]A�`�=P'	L�|�ZDhV$��s�}�3�͒K���.H�͇���L��ؾ5B�!���<;Y�{ROM�*R1|�Te�֕�M
 ÔjW��p������"`��e!J��ΪgC��=eM*�0!���:1�^��P{��5��a.'�5�u#�W[BS)H��G����4��j	h���|-�N1�@�����d���b�[�ka�,C8�R��ݵ��VD$��]�O���8��l�.9��R$�I�dG�0iV�\��Z)��M�Xd1[
��Q$� �\8J�4�V���*� �� #FZ���OJb/��@���	G��*8��H��9����1�XЙNxT�O�Ƌ��:��E�ML傴��p3P�p�[�(6����2CQ�䉍h;c"���e�T�R���̫"��Rv��X*IA14-�jn,����j5�KL+0�Q�J�kH�����h��$e�L-h1R*b�(�n���;k�ܬ�e���k4+��m��rE8P��_��