BZh91AY&SY�[;� ߀Px����������P��]Q��8cjd%A(�*y'�6�l��C@2h h ��di �     ���j�b�У������4� ���0L@0	�h�h`b`�$&�S���<M	���F�� �M�ҾI+�D��#&1!^?�⫚�/lA��I�,!2��)���`�в��G{UDa ��G��:|��t��.y�t��"��E��'gRK�+œ �"�G�{�N<3y\/f���>��9��۷622br�Z먠q:-������	b��V�)Z����3��/q	d6��yD��鶩���M>O|��I��*((����C�Cu_BE4ExuU�c���9w)�\̓���x��.�W.]f�25x/�T��� h����	-���������aa07�SK��X�E��̒`@�H*�$M�0��P'+�7�&�vX�^�%�aA�B<��IbeiP�����>2��)M�K���ZsI���ʵn�ԇ!�HZ���I�%�ST4l-��(��Ace����h�� 0��(�`�=��{��r���6�m!Bk���B��#�
Bw�j%J$��Xcd���hz�/"&F���� ���j�d�)#�eZ�iH!lҠ�a�5|��Ch�������>�x3�ow���A�7M/���U1FE���9��'>'�#Y�)<Ϛ	2�B��x�1*�N���2���уp�z�_��a����s�xvM^��oqړ?�H��hX�iz�ᖭ�����a�ώ����=�e�I��iT��D�F�d��a�f�gՄ��)jmyf=����~�%l��٥��fƅ�;|z����ȉs�mrj�L��Bb94�+�C���*�eW��y�!����&�����m4!�'a���=�� Z�l
�ʑ�p@~�8|�&�8A0`�b�|��G>1����e�rіҴj���&��ж�2_	#&Q�pR?�Z�&�(�&�ȥ�U��O,�*�͛6�����I�z'����GKJ���p8�F�+p^�`���x���p���p��Y6�
:��"���XtHF%���Xg�f���`�Tf;ؒZ�ZŴ��C��%e��OC��ڐ��|~��O�ɱ�k��{79gl7�77�y̕�����+�J�d��R�N��e�/n�L]OC9Й�َ-Ci�9r*cK��"��o��(��n�[���h���r�-����ޒ����Y���iT�]��t����9uh^g�h]�޵58Ye@�����i����i5'z�L�*���1n��l�,��Ƿ�MT�r�1�?�N5Cj���������"�(Hb-���