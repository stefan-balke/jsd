BZh91AY&SYp��& e߀Px����������`?�Π  	D���Q�&�zL�C���#�2bh�Phh	��@44�@@  4 q�&LF& L�&@F �*~�Jz�  ��    q�&LF& L�&@F �"@�b�=@ɩ��� �	���=��$�%`���G#b�U�Hi)�$��_��pxM W�
ɖah�jNDBh����tsc�,zz��'��mۇ9��~j�S��kZ|�`�b/'?� pp,��� }���$���ýEnnݴ�h4�r��+�n��8p�fS*2���Α�Q��F�<�O"st|X�eN����hB���ЅP����!�����[���r<��.� h�A�zOd�m$찜��d����T�@JrJ
dn0�����	�P��]� m��Ѣ��4�[ܕTAA� 8=�'$��I�MZ�$�b1
�(�B�8�鉫!��Ҧ9�3�>V�U�.#B��X\�Њ���AB�Qt�*��PSo��+LWh���3�wC�B4 �B�D<0*�J�r�<@�t��F� h�)��yeey�)�I�i|#��	$�Z��a��Sy��a�.��,m��#Cf���`b���̻Բ�b!g!_9IV���+/k��7� �AUZ	J]��p3�����$Ȼ$LIZ�0�(�j�$�����#	i%D�ilM&���(��(SY*4��_M+{$�����@QUH�)c^U������CU�K�s��k���:�z��>6h#�����1�0�`����EfS}����fD�N4���u�?4��p�{�{�T�p�d�b��@1��i̯��oC�2@���	�Ҿ#3�Iw"�^� ��f|hI�ׄ����}*��A��ʒx�%Z�~J�w07���f���DP��-��-��L�0�j�V�2=L箴8��.0W� �CBq�C�xX+��A�0�\d�(
�=���)�s��͌��G-���_0g�H��uCF��7۟��`���g(3W��_ȶ�������{A �:�fǶ��<8�łƐ [�!��w ��S�~'(�΀���P``L �'# �7<f�-D#�%$ t��" ���<d��P���]!��N�&����H"l��ǵ^4'�>fhA�9�@=��@�>�U����DѤ�c;�/l�������a�$$�Rh�a�wq!A"`3钼��x˃�WuT/�N���$1���(�Lx�hPf|4�U�V��R14���MI߫��T�!�C8����5�\�J�_bAk��,0�MY��m��f2��#w��i���z�9:�����	8��k,�l�� =�lmx*Z�~��fB0hZ���H�
�$�