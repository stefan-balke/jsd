BZh91AY&SY��R� $_�Px���������Py������%Se'�CD���d=M�C&�h�&��$        ��S���F��Q��  ���A�ɓ&F�L�LE F���S�OG�<��6�F@�̲�P�t��$A����DA��	��r�q��a!�sd���M��ґ � n=��Z���|Ol��eT�&���^��o=�����1�:�`D��/c�����&�Ä���3!�X_q��1�Q�"NZ�S+��b�<�@
�,��
����[��� ��
,!����!�&kz\�o=���S_�zi���Y�(�V�[�����g��G;P��5@�b]nS�')�,�LK	9%��
8���Y��&B�Gp��n��ҝJI+�T���Rb!@QV��a��XFb�B�[�ȽU�X�nI��K�
?����7�m��СN��ZK��G�;�J�IjvX��1��± P�'r�6�6F�Q!���#��l�PP0�l3}&hH�ojV5wffXT������2e
h�v��M6o�h�X�}��-�+�Mq�+Y	f�}hzH�����V�e��
�M�F���r���p�gxcD�A~�����f���A�A1�^w�K��)��APM��nBe'6�"�	�cUP�hD�{;��KԒx�aR�R��wZfR
�A#��qjbd�Vi��"���V2�<��ѥ��25,�$�i8^M�
�:���P�Xf�(���C�K��g㓎ЮB��~JB6�u�\*��Fh[CcÌ�)JG�����B�����u���� �C�_��JS�mPтŠ[����x ��S�>����a�B"cAC%9��`ܲ�a�$�b����"���萍/i.�p�+o�r�BH�EĠ�$��k��	�x.㒐��qH��y�ʡ�bj`����d������2��q�*E	�!Za��PY��3ᚴ���-�s�Yy�Pm;�3�#"1�W��$<E��ؘ�V؊�E-�YV%IP$��0T.�dS�^5SU��!Z�\��@�2*�(�iy���D<�փ�]	�ʥ�QJ.�5ݕU>��C�K��
�FS�.�p�!�8�n