BZh91AY&SY�?�L P߀Px����������`�����84i��	D�M'�=�i��!��z�h4�h5=4RL�h3Ԁ�� �0`��`ѐ��&��B$��jd�z�H4�  =0`��`ѐ��&��D� F@Д��j�	�<�A���o��Ԓ	BA� @�r{�F�� ɡP�$&S\���p[��
���@&�֤�D ��_W8t��]�>�������s���6���71>fc��t����gu�+D �ǥ��z��nkA�B�IG�M��3��=��a�����˨5s��l;�`���~Ya�u_�Arj��^`�RFʡ�;�fX����'fk'0�,3�B70��'"RRe~_*����V��	�v��|��@������x'�/�0HN��; L�����v|et�f����9s򖌞�\Mo�mp�_TMo�2��(��(���` ������Z�)5���m�R���Dڸ�&r1WDm�3�ӻ�dQ���"�0cn�M^|A	�1rwŲ,W&�MB��T�ik�M&x�8mC�f���Sjq��fBړИ}�".7m�4�S	�Td�e��D�S��!M3�-���Ն�qS=���e���������eF�y�/�f�l�C*5�mJmY ���\5�4��6�>m��2��}N��eLM�{r,DV���w��U3Y���F@�I�]0�Њ'zȍH27��9�6m5�lc{��CI
㳥�j���RC��T�K�8�i�lm6fj2Ӑ�u+��C�H�e��.��L�F���bcm�5SM���X���/*((F��R�UUEQ%Ю�W���_�i~I��Q��iH�~�/j*�p�!�nsZG�EA��Ɖg
}��x�E#��^L�KU���mj�g��&��.&0QJ��F�$���q�r��]�xc ����bB�B@b�ڈ���6�L2B�w�U����rK�	�<D��#k<�Hd�Pd���d���f�ҁ��dyv$�	R�[�F�	NzK�ڃS!3�����0F� Ԛek��EYΰC�7���^Efuoh��m��1$��P�,
���{m���J��(K�����U�@1!t����T�$���ur��׸$A�hh�\I� �ြ�tj\4�v���$ա�b �u��P�^����)�݈`gXN�Ӑ��:��8�?��T�Ӥ3���D�r�KvpQ�߷�� 4k�PE�x�c�B0^�Q��p�gL���T&)4P=e`%2 "���$'�zD��0���xD4�@瘭3!ea�!��`o�}A�hL��td�B| ��p@��̄��M"���\Xs&XEg*���i�:7��ƃ��1�y�Xm���k�~qRKC}�`o�EeT
���t�2f�1�/�I���}-��WX�:���璢��F?r���^c�ybli4/܋փbD�͊‰� ݮۺ�ב�N������j4+���H�
���