BZh91AY&SYn�� k߀Px����������P~�M���6�����"`FI��Q��OS@ �h�i��i(    2d   HH@��bmO�M�Hަ��P �ш0� �`�2��*IM���I�ɢl�MdhhF���h�`%wH��#��W_��VL��b4*L�S^�m� �Y h4,�&��#����n�Sxn6j�^�_��^=��-4������ʙD����q���+l�t����-�ٚiwR����p��6h��K��Ǯ�ɦ���2��Ŧ׷2�v��DI
u]M���c�Y��������ndyz���(�h��v63�����Ϫ�1�&�-J��:�M).��AC�u��r�+����d�֭�d-�a�"Y��՘��͕ya�bv,�Rn˝�\��x��0�
�B��gz� �	2H�v�-��W�2�t�VShR)Ud��V�P��l� �VHh�X�Z�������W/�dk�\6˗r����R�9���lc|m���;l{���B�ȎT)�R�,�k��xv��a�����2 �䳃�&)�EP�T5j����PP0�u�>�@1�ѳ�ͩ���^x�g�F�����!���7a�I��X�s���$��j4wl:��S��h�w8�M�_!#��&%�pG�5���O���z΄��T��Z;F㚵=Zs�K���g9���Y2���ތ/�m���I���H~cz�����N
g�JR����}���=F|�O��X�z\�m���ټ��y��ɭn��ˠ�݉�"5��1J`�Y�!��ό��-9A��m�4':K�za-�o�m5b�����<�j/���Hl�v�S	�d�,c��/I�C��#$�T+�P�n\t�-!j��"l3wۈW�O=�UX�0������l%)]�$0�WP�}*\�qQ�~���Ƌ���u��+)u� ������7G�{H�
��	�PX��v��%�.�a�>�8:����*1:X�[
ZŶ�;n����$9\L7Y�eH�y<���֙�,5�X���n�|8+��*%2�t;�,�V�ڊ���kso�oF�陋���6%6�򙳗FӺo���e�WL�����ꛗ��o�WR&���A�Td[eOM|%��;�c'j(r)�dsY����I���;�"���y�$�zG5m1
�H�3%����Ջ�N�ّ�p*':z��d^~�w$S�	��A 