BZh91AY&SYX�oE +_�Px����������P>�ɚ��bb�D���1L)����z�OS�� �1A��4�����    � !"j
z�@i�=L�Q��  ��9�#� �&���0F&
�M0&�M5=2����@���Ҽ�q�E�&1ЖB���ج���2hT0Ve5���0���	�`�#{(4qN�cm��L���r���f�d��/!����X��B�$���2"[�++í��5��]�Ԭ�L����:�����0b.��6�Y�沀@��u�"PV���\�O��D��zV�&L5�����T�����[�j/J��\��\5�ƹ�.Ŗ�=��ΦF��#�,�bk3�T�@&kD2Q&����Y��Pa�$���Lb��e٢�#$7ɘ������3)eC5L09��f��ÑM��������E�3V��m ��#cަ�m��������P�vH�B��9(�(��ȑ�����c*��o�.�%AG�HGيH�eZ�g��E��K�lbLȓv<����~5����ۻ8o���tt�r��8���y���Ĭ쮒Av`�}gW�*EnS����f�����Z���I>�wn��w�����
c֤��hX�iz+��N��R�Ф�q��~���?�3p�yv���Q�Nw��My�a��23��n��C��ԓ�p���k��4F�Ž��5DK�4WU����4u��+X�h��*Ȟ&k�JͰ��g�4�m�^nc1�z�Fº97����c3%�ޓ��1�}��$���v��9Gg^^�>���o��,�!�dT.r�P1ovMX��һ�d0�nE�	���]������ݣ�������@����;F�/�ZlA�)aF��Cj��Kݸ��W�ؼI�ac^�r�<�,HHF/I�!Y$dB��*d�ݒ�j��Ak��-������ޓ��\S[�Z>��G��Ns���k,6�>l=
x�<0Wy�Q)�c����I]CYQ�R��Ot�L"�-�����g:�?fF�T�x����գ[���n�ss�ΙZ2�p���e�/0�MX�ɣ�Z���SQ�R��dp�ɣ���2���-1�R��P�2D���f,�%���/F&(���H�Y��4ip�LˬУU62�à�`d+r���]��BAc�