BZh91AY&SY�m� n߀Px���������P}��5A�2
(E&jb<�jmM4hi�z��hd���A�@ ѓF�h� ! �!��zSF��� ����(         *�M!2zOBeLѢyG��4�� h�M<��Bd�$4 tOBL��bc���y�T���J�&}�DF��1�e�����jD#�����ǯ�=�>�c�93��vv�Q=}�õ��h���ukP�j�Ͼ� X���No����mћ�q�v��R#`�(akX*Z�j�Dۈ�-#���@�N���,��`g��P�ײ�/�}���� �AE�N��vB$��ӹ$Q�I��#ޛ#FI�S�X����Q�k�&�S8�=A��2���8Z�wF��X���jʼδ��P�f��Py�`��'��0c(�FF�JS;��q�Y�sgk6@���U���gR^�J���`�Q:©'aKpp��%Q2��a����[R7���O�lcc��m�4!����@|T��"8���(�(����ʰ�?�,Z�.21�k2�)�䍔��e���"Ҋ
��g�`1�l6g�ڛ�~��ݏvx�����!���;�m2K@��,Y���CmJ�Z@�f������E����++)d�p�jL���yhr��<�}�����>��N䇸�6�ݳ��͹8�*?�����������.���[�.7G±�"T�m�LOgt�����|
��4�Ȗ���:�({L��\��-\\�a֚Hg`�Z��*�>fv�d83��d��J!�0�.u�F%�T�9<4�6�2�"�
�=G��aeP�y,f�z�+���~�F}+(��L/l!�n[�+�(��Yȗ7�>�����n:�9��
sG�f��{߳��L5�ɄGE����	��~��fL�5:�knMq��#%�y��t�Ͷڴ�h��j
yz"�TX��%�	�}��H�j�:Fn��Ф��z�)iI:��w(D��0�<����ѲT��[��=���G��Y���d�d�N��%~�[���'�	�����w�E�&���������qsx`m;�gW�2�1a�P�m�:L��:�zB��:����Z墳�W&v�Ĩf��d� ���:1�#�¹9ʫx(Zѕ}q^وs�ηv���=j:�˚dnb�ij^�
:x����3�0����L��F�n�8��H�
�� 