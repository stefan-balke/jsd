BZh91AY&SY�]� 8߀Px����������`�B(u-.l  M6��a � �   5O	�Jh@h�i�@@� hh0`��`ѐ��&��S!�6�e=&�����zA����&�s F	�0M`�L$H!d���)��4�=	� &��u0�A ( ����E��hR���I���M����e�! �ũI� ,��s�:9���]�Gι��e+KKK+K�	<��z��(��9}��X��_h ��R�$����1�m����I��i/� ��<���vL���A�L_���Ñr�9�#+�0��{�bHE���J��A�!r
�$��7�"4L��9I���[�����RB`ǅ��uR�ǝ�宧)U��}(��.b��92�lI+��R����2�}�4g~���A[0��2�G=U���p1��h��V�#�ʒ��9&`5s';�)�i�njX篇j0슬�j���+&I�&�����-T���XƖ�ЉU8$��!܏eP��Y��e����!H�m1H�lf!Vs�����ƭ]�0\[�Z�Ȍ+��0A_E �A�rp���I�2w����S-��ɋ��*��gSC;��2�q*!�(�!	�E`<����Y݀ Lʳ��ֆP,*�z�C���r��
�:5Zq�L��ң{E�:��;BB���C� 왗�!}�Hq($�;~	���e�L��{���M�dȆdbQm��H�0p4f��)�.�Hj��.�J	� �HC\���c*"R��:�KNH���������y, _��':�6�"J�m���{&h���������&�#��w��uS��9�O�CB��!2���d	����ػ:���zċ}HG�� �qq߮�B�lB���Լ�kڒ��Q=��#�*f���%b!���C��� �-�xP%Z�v%A�m;Z�uf��A����њ[���%��nM 2\0k4R��P����·>]��w�0�JA`W�>�0��a���4�
AR\Opz��=*�#���Ldנ�8X����-ĈtGA�YJ�d���QT0S^�g037�~���֐��^�1"�>u��Ǧ���!�B\�ݴ�G�#�r��@���m@P`h0����V�w��`� $p��W����;�,6	�9L���N�&��ib"l��l�%�؄�S�!&���H04P4�>��C߁�Ј���F�j=H\����CPЮ ���8��!��ќ�A�䐍!4"g�J���G��9�q�`f�N��x�h]�4�"c��#Ѹ�̹w�a��$���a:�ԝٸHEL�3"���5�[����XH,�hGSt�"�XMN�
!���O�H����ɤ�G��oI�.h2B$Xe6f*$a$A�(����NUK,���N �0hY���H�
ˢ8�