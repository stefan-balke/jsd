BZh91AY&SY�l� �߀Px���������P����C84	 a*hD�MM��L	�L�d��Ɉɦ��OBb*        M&D@Oh�ЌM3S&Lsbh0�2d��`�i���!�*IL��2d�4�����6�hh4��h_	\"%�C	��Y
����]ʪ��`�S_3�p����г�GCUD�$g h�s��8��|��3�|�G��c5��O�k��7�Y�`�ݹ+�U�+�(�8�UK��8��'<�{�pL͇Pwڛv��;7Sx��Y�����tt��Ea|D���z􉉑=ÚX�̳f�h�C��� ����:L�y��ʫE�l�]^�,�f�k���E<�:��7<�p���cLA�aBgxa�2glҫI��?ؠ�/S�����l;Ѡ3�A�PR�-bJ�M���Ro`�)&��)�,$."-n��km��UpQ�-�!�Uʄ$��c���M�aw��SL��Z鮘�
P#��Y�ib�`�RpnA�����61���m��tw�_ x�/'9�P����*Q%�ٓk�����#Čm�(�$`UU1�H�2�FX��PP0�p���hCa��3u"s�\�C1
O�L�845����Ir?IkILq�T��u��F�K&�o(*!��/����rcX�jN�M����;./Z#�8y7�N����>y��#�-���lѱ/;�.�sbɯ�ϖ�{Yu���S����H����N����K�����}T��{.�%i��rͨb�H���heRʹ�`�˞�52̄oLV��0���b.r�+���̚g'rZ*��U��t�21�+�����s35��������a�\���\m];Gc�ˏy�oC�`�ϔTcu�9�����o5K������Ӹ���m���#��m�,[D��gV�q�ѿtb�z�f���7A�H��cخڣ�;�l��wb��y��_{h�n��S����@ Q���� �ĲBB4�i2H�4
�;#3�0Z#F��E��Ѭiz�"V۶���i}d�)+�y[������v���X��^sb�S�[�����Q�R�_F�5���������f:���Ľ��T��T�J_Z�V��h�nTۻ���юs�q��+�/ľ]\���#{�,lr�SB�����\��d�y�]����u��a�R5|�~�ꒉ���m9=KȽ��he"�j�8q��㢪|��T9�R�:3�(?�ܑN$-�=ƀ