BZh91AY&SYJ�9 �_�Px���������P�:I   �U4F#� h h 2   ���a2dɑ��4�# C ��5LңOS�OI���S� ��d�A�ɓ&F�L�LD�y
bz��L  4�S'��M	�@�IJ�Ͽ���Uj!��0 �M��n�1"����JPȄ��ˤ�W&�|���P�2��zKV���Aegi��O.=:]_���{Ǘ9�f6�EFX��sy�#�[u��"�2�����lz�j�u( �-{n�'?�"��xl�;�
`!%W��k��.#~g;Gs[*a����̽VV{`�vEb�A�D9'�jא�:.Ó4�:��(Md(d�JE�Z�I^�Vjw��5�T�Q����V�ub1�pЕ���z+��s%������I(��j���ψi�$>i��X�*$bQ�K���ViE�D�J �Ciaye�$��k��Ƀ6+�~�$�?��_Yu�aٴ����-up��V��**'�Pi�Ͷp�唄�+��w�4aIu0@6��¢"���XB��'�zږ�������`@lN��6�SH2i�5�n�_Q�ޒ�¥�X(����P�Ѣ&s&��!Q�b���dw��I=L�J���1va�}�l��&B(K˄qj��i�m
q�e[B���^��WjC����A��h��m(td
����|/��m.26��Ab]Ǩ?��6&�9�]d��eQ���!M��YBG5��YM��y��*�
)��7�0�t�24}K�z����Rɢ4��@�ר����CKR�!W���p:J����@����%�T`j&Z9���5�Q��HĀ $t�P"A2J�Ȃ ��̅D��*�1��9�&�h�z���� #��7�=����0���A!������dh��1��o �4&z:G �$��h޺�y��&(xlX����WyjӚq�H�aG��f�q����p�*�+�p���X�BjN�8��P@ͦ��1�`�eC�K���Z����0�Tv�u��>/=&M&����m��E����$A����[_#5K^_�"��(#*9q����)��Vy�