BZh91AY&SY��Z  ߀Px���������`�y�nÀA�4d�(��O(�OiOPѠh4�@� 	S	����@     9�14L�2da0M4����$" �"4��'��M  h0�9�14L�2da0M4����$� &�i�@�ф���z�@ i�4�BW��D/ ʞ�)	�
���:8����-
�$ZMO��8�HKa���@�+T��@��w�/G����OO��s�}m��l�&�l�Z�kKr�V�zU2����av�ה޺���)�lm���ӛ��T!�Ȃ��r��5����:#�'1�ִ�fFhY�;�7!�;�Q�_D.)�>5��ގ)��V���Ug��`l�3�c�<ȭmVU'��0"Q����LATPQt�:Y�8��nt�/j��}l�;�e�F���H�76Mf���:�M�	R$�qs���kUd%�+Xo�9-�"����dlyCZ�7t=�5iSF�[z4�-�0���UNlS��y�DL����{�Q4����*��*�̕V�e�Ept԰���4*�E��a���3ޟ��,�$`Ѝ�+c�v��=B�K�6�9Ѵ�@�$�|ap�k�d�Y��a�&�Pt&"��ȹ�Iz�M��²�ɩ-�"��d�����#����~�o��ۊ�[+��z��3��;`��dH,�|=��ֆ�w��s�����mI���u��Iy�9J�x�Z%J$�� �A�8S)�/B�rz�RkB:LM56�X��4Ӧ� ���m�(^�PP0�w.�bI�P�Wކ�����!S>+������xzV��a>7J�k��>#@h�S�g�9�>��cʳ����e�ҁ���}�;��U��ER=�}���k��>xg�TH��B�&�f+\�mյ/7�5����$���W��mrO.șR~�W�$yG7�W��8P�?̷i���}>fB�O�$��+9�^���bK�u��{��Z���+;�XI3H��L�`׸p����FW���8�����s?�,�TT�Im���S�}cY\���˒�잷��?k��QQ#���rn�C��~�FZ�Ba��AP{\�Z�6�L���+��4y�r~L�x�m���:-�<���aͿtq�S]"L�o�6v��GC�z����G�`�CJ��V������X$� (���"��<f�D�`�0���2[c=���tZ����-u(�����[vqĎ�����Y��2)y<s�\�qa��{K��ή�b�S���:��"���TT�YGWv葉�t��X��K���N��ڋ�R�B���dR�aZ�$\�R[��z�ws�,�g`�#��h^B�=��BFM�prgB�Qa��]�(4�i/!���SQ����.����ZjJ��gCi���IQ�ַ2M���σk�v,i����TTL������ܑN$:~�V�