BZh91AY&SY)��� 5߀Px����������P��d���2kM4I=G�O54� 4�@ ���
Hh2d �@�4 j$&���MOI�&�z���40G�F�c�0L@0	�h�h`ba"Bh#!=)��O$�z��OP2h �6�$�IP!2�&�!D�_�l�����	c �$Kg��� 【�`�2�!GV��D$����^�t�<��C��M�kv�kgZ�������yw�P�pJ`���m���[e\4�f���h]e�g�Z;=m��?��ʌ�i��a���1�d��R(����O�V���4
ݍ��HUD~�r���j�]jg����v,���NrH��oι��@��M�X	��w�+ԑը�l�E�0�9]Ѐ�h���N��D�ʣ]ЭZ�o3���3Ja/*Dђ�l���/`fTV�Å�[�.��0����wL��z��T��� R*��:���a�×YZ!��#0�@paD�Q@9$:A$��s�'��0ڭ�����TQXJ��v�qu��eD#��s�t��勨g[}��5[6a�L��%�V���҂j�M���1�?Q�(�"�UV�QGN��;�N����,��t�WVUbȟ֯<[T���b�@h����SЪ`�ȪALڲ�B}ic)r�ke��Ϝ��Xox�ֿ=ywg�nӆ�)ь!�>����� K���YX~g����P��y��yb�,�n���8\�Jr����q>�<�͊~8�)%��zu]}��G�;$[�bK� pP�e��d�� �9��WL"6ց��Ip��D
��!�b��u�0�R%')��y�Ԣ�&�G�AvYu�+�F���Ppd"(x_-��Q-HL�!�)d.��K�Ί��g�Ҧ�wXM��c8ȡ� �Y�� ���3���A@XK������PIt�C62j@�ʨ���;�>rd��CF�M7��%i�1J�LD`%���߆�uLX$��V�p5K�����w؆�x����$�a8�hԧ�~�(�a������`P�li��Y�����y @H�%$(r�eQL���2��5a;f�.11�AI���* D�����P��ė������'�w.r#$��@�:NZp���i��;���:�B��I��fs=<D�ࠉ�[��O�-��@�`�,w�N�̉b'�0G��J�d<v{��A����VB,�5��k"��	�;��PIX_""&�``5�Zl-������h��x�0R���P���ש�0,���I�f�DH��,H�H�L�=�`���J��ś�� �4,6���H�
10�