BZh91AY&SY��"� x߀Px����������`_ض�a�`P( 5SG�i�M�4� �`�C4i* M4 ��0`��`ѐ��&��S�DG���=A�A��  s F	�0M`�L$H!14�# �&�z� �h�^L=���T��H����G#M���Z��HI���M��Z4�XX�GKRrDBd@\���[��3���m�����e]j4�ͦ֗YQ�m�����@����Z%MP����s���Sb�塴�pܥ�����x2��"�,-2���$\��/�AL�iC�2[%73�+C��hB
�d�%PЃp�*��Ag_wθ���غ�a7�'���5��[�hM6M�ƩQ�>�P��H��n@���k��u�΅�@��gu8����l��br�8Y�B���a%����@�(@�Ebτ��-����iZ�N��
(F2���BS;�9pAj,F��F2�T02&��հ�P*>i@�J�H*��=.L]�@CNuGL�u��>dh6Q[9J��-BܒX�$��p@j�w-�
<iX�]H�4�na����<�KK3�k��F\�H;[.��a���*�6�W �e�l���uA �"説@I'��֢7m%����SD��tUF�8�LKڨ�a�%�"�kX����%�Y�I%&Qn�v�%�.T�u%����B��	$����R~?춿�3��i=}�3*w~"�i�p� �!+��|�Y��@�����x�/�>�l��$I�v�g$P�8x��H �y�o�y�Aq���:���@�1�`^z��q�׆�T9M��H�	�^W���W�͛�S�I��	�FL�xP(�9�}�M����j&h��� �3u$�T	V���Lv�_3Y��`Z��˃T�50��	�����JTs3���'�a��oq"�**�@�e㯨18G�p|�k�Jb��.��=��2�KI ����F2k�I,G?���׸�]�|������QmT�a3�37�:���f��5$�Z��|����Ek\�v!��� ��H�Q�G���9@j�\s%��P`bL0hS��V�3��L@�(G��X��6&I`�a7�.�`�"Lh[TN�&����"l��ے][P��iHszS��0@Hi^�����Ȁ=ǣ��3i�����#BgW1�8���8������j@dq$T�ү.:��Zy�����N��8��i�"1�2JCZ7�c5�w[�VB,�/K#��,'P���7�S4�"�x�
MbP8UYu�����Kd�TH(�˵O��e���li1.��氹��	�,6I���g� ݲ������U�ۿ�d4�
�K�w$S�		ߢ+�