BZh91AY&SYL��s @߀Px����������P>s���aΡJ�@	$)�M�I䆙4��  @T��(�       	LRi51F�G�4�� h�@4�& �4d40	�10� A54�?%7��
z z����=����H��!TB P ~^��r4�*Ф�%1&I��xͷ�0J�X���U�[	Y>�٩iզ��}�����D߱рk��X�ꖑG �{���H�^�}�f�dgH���1"^(��X��[�ФS�Rt)��܃%��w�Hk�Ԡ!X.�ⷳY��+w�X�\���Lspc6D���E~�
�#iF,�-�'X�����Y
1fYL�h�(��S��)KG�#�B��)����4J*��ae2t(��)!T��Pd�*�Je�]i�&I���"4��4�HD�qTJM$ԹTbx3�s�H�j��/ՙ*�@��R���&c�|�$!!	hI$�
���-��|<P�_ ӌ�K჎�V:o�"�J'"��H��
15Nʨ؈"�a�e����g]�E	Q�:t/����_�K$�nRw�
F x�/j7��ǎV��!��Q!�-��p����/�n�v�=�3Y���;�It����� � ��#�A�1>g�5c�P	������8W��qN�X��Ě�/���K��(7u
����d��j��T;����Na�����4�:��Р��ESsTI��1jhPp0i��XR�G��UqC��y2W����q��tf
�@N]�0���P�	��K?��(L%�A���$���\+���L�Ψh������aE�2S>�f�f��>e�i�f%��6���0�5�r���vHW�K�)�F�vG��K:ȱ�D�C���+	a�h󖢫h!�ܦQ�����D��*�hʎs*M�P� �� 16�ܻ�D'���t��ǯ _�1�?��(r�0A�d�c��Pޜ��m!1N'Q�,I$�@d&� �;6	i	�ɞ�U厓��p�*����s@�7�&@4Q�$9�0v���3ٺ�V\v��"��Rwἠ�L$8n�д#P�i@�@����4��P�� $����i|^�[I�w�p�s��IH��l��M6m����{k�اk�vs��A�`а�#�
���H�
	���`