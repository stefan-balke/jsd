BZh91AY&SY���� o_�Px����������Px�u�08�M �F���	�2z��h��� S@���S�@h     !(�5=Bh3Bhɠ�4 ��9�#� �&���0F&$&�S�)�?Ry2z��z@ hѵ6����Q$�� �!A�������f�p)��~.mæ�%�hX!�0�����HЌ$�|�ӵ��}�/�I~l�JjX
�蠈_�m)�K� 6�V�h�D2�7̬D�8O����	�D���8A!1xCz�ә��MH��#�mI�1Z��9�!WJX��G�VQ{@�!t2�L??��Qŝ��xq�ߤ<d��[e�%}����d��qE5T���+��,��n�eLA���M��s"G)Q���]��	J�j��p�\+Q�;x	��B�����V4�H�dU\0��<� �T԰�C̑e�v�8�C���@#*�%�/4F�C���8Aas�֨1��g����{m���u�N=F����7�m����5�g�;�-\�r�@;�5�QW��B�ܱ��ƓWHܐlc��ܑ��Ư�)B�#Yo-���Z�t���9�6��n-���Wφc9�1ɛ,xa*n�O��	�	'����z��;s��VZZ�F��Ug�3������m����[b�^��HHn�gٳF�P6�!Lb����	�Ծ#3ޒ��� ���ə��R�	m`CG�s-i2��T=���ojI�@�km�Tg/AyV�͐���t�5@@[S\����������CN���p�+G �M���E���+�? 4��va���LP%�x��O% �:9P͌&�$���u�W�g���ф�����iE�1S^$� ����0�K)�R��ʕ*�-����a(���(�Dɍ,��J�BY� ��=@4t��=P�Aa�A��0��NfAXnzf�I+���PX����D�h=Ľ"�%Vm,��9�Ԡ��P�X �� #�W�Ի�!<���Li1B��<��^��&��`��������=� �hL�Q�q	 ̅�W�:OV��`L�d�,9Ah`/���hs@Ύ#$1���1�2����͛��U�V��z�p�E��\	��q*a��A�H��4@����Z��\H,�`u�I]�KAbF_Z�sH��ݤ��b2<�7����a���2D��{7`��U,��k=f�f0hXb]���"�(H_�D� 