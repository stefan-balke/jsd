BZh91AY&SY��A� �_�Py���������P�71�r�@jh��SM=&� h �  h Й ��    Ji�"i6�b�     2d�b`ɂd ф``$��D�A��j�=M����4OIy4$�%	!I"�~-	H@�|Q���hRH&���_߉Hn�bAp�Uab8�&�d@\��}8uj�V�)���A���t�Uް1 �ھ,V�s��J�4���Z�U���P�x�_��8���Õ����;3$�x[�ԭô�oJd�~�O��;��I%e�����B8&0,�k�Cpܷ���\s
��`Ǖ����r�p���%�n�5�@�B��˕h��U�l풢2���nl7*11���B�h<Hz�BW	*�jڀ�-S3xVtH�Q^\�^���E(4�'���t*p^�JM6fb�7�%|4]FA|���ʮ��j�NO7x��B���&N�P�2`t
ı��X 9;���4E\��(	��9&Z�o[+eh4O1#F��m�ָ���;��c�v�m��PA����=rK���.F�=�K�LӛX��
$)�'H�u�R�̤M2fD<`�$$$L��PGMC�n	+7%GH�rQ� ��Bv�E�9�TLL���P �3-z�Ĭ�`@�u/Mq�1mx(B���r@nE�zL����6�{��I��|_���(Pk1&\�yCvZ�+���r? �P�s��!!��f#�?�^��*A�Al��Yg�z�3���%�^�0�(���ΡQ3s��d��f�E��� �O�$��%Z�m?ƴ!�0X��{۵�52B\9���eCH�M$3�D���JQ�7�z��Z`�w6���J#�PX���v��ZhS	w���SF������I(D�/9$tX�6���n�^EF��!N�[M���n�U�iS<	�`�o���}嚴^ku]zš@@F��9����V�hΰhA�v��: 4u��?Ca�1�ʑ�*����Nf��7<'�S�-��8�� aD�ס2d�zIe���G�
�.T��wK�(�"/6\iG�OUqp2D�fՂC�����\g0/Dë�#Y��]���B���Q�2I \�t��&���:} V�L�Ү,;9hu��*�ׅFӢe��e^4P~Fp0���ճ-�"��,��ed�	�&����PS4�3Iz�9��⁕e֒,.�
(���S��10�=�i1/�p����f��P�� fͲ[mmx�,���A���\��U��.�p�!�n��