BZh91AY&SY�hOk ^_�Px����������P~�h�eld.��QSҞ�=$=F@�1�  �A��#G���h Q��  ��T�F�A7�SMOI�m A�C s F	�0M`�L$�MaML�M6)�6��4 �c)�tEp�ZI%�C	�W���V&r|l�
��`S_ؿ�6��hY�=U4�2�����wI���8ygO�m{�6��ڙD�|}�\��۠�r;:cn�yNW�|2'��o�vq�.�E*b��[M%Ŀ �E��n�S���D/��"X2'�R��Ȫ]���nω�wa8�J)Y}�M��}�Y�M�S�F��hz+A��b������1�
�U-=��s�a@<�
U4��`�!^x`,)�)\�������N�8���LJ��U��A�)�*��g�JZeB߱qµ[�%�2���L��V(3Ir�GS�`�z�*���+���_f�g�N��x���7��m�4!�c���.��9P�;��%J$�����ָY�0Th��$nH6VeF��F�:ڰ�a���#]n�DQQTI��U������J�sU9�W��k�=�� �]h��}�%>%y �x!n��S��8[�W�,�V5�\*u��
�l.P�SEIV���b��re�P��c3��۷>ļ��u1.�!�Y���y�Sw	'Yy=a�t��^_%9�n��S��6<q���Yg�'\��V1Ŧ�i�1s|��-C�ȉs�eoj�e��7��]5�_V	��1����h�z��UJE[R��a��Ԯ��v�S��XP.Wa�/}��� ��煌��)
^���;CFr
�"	�7�%�H�W:
ryh�f���ա�2f��%��]&�x�3+^cӻ,Rg�/�'2�w���u��k���X�l���40-̗�h\g�.���j�n��)$�sꠊw͇D�i~'�a#�-�|F`ݬ��⦌L���X�����+o.��8
ih��Ĵ�.�쇳Kt�n�6��F�K�e��lTJa��t1A�[�kJ��(���˒玹�����2��-y�9yU+���QC��E��7k�s���g�X�Ɓ�Cx�g,R�Du��R\aXca�!��5�.�gL�����際��2��W|���j����J�9���j����&�Qg>�w>j���/���5*K��@��ܑN$"���