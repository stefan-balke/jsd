BZh91AY&SY�BU� �_�Px���������P���jN�� %xj����!���C#LFF h24L����� ���  "�i��F��0��  M sbh0�2d��`�i���!�*I4D��O&��yOf��  <���+���F)#2!_������\�0��� �.I��I�7a�rXhUU�!���rEb�nË�?g�s1�_ln�c��e��1�	d�ׯ�E�����Av�1Lԑ��CI���Sps1��M��j��g6���1��!X�6٠nq/�QO�C���d�Z�+�IZvsat����o�(a\3cqq���v����$4��=Q�<]P�+���ݣ���
h�r�/�A��ڧ���.ˮ��fm �a	ޚX���ږ�4��C��V�a�Ba$N�q��D'v�
�Ţ�^�l�)8"�øuN&���D���..���b����OBJ�U�2rMi!5�vH�EPWEU2�y�k��KhE����z�������j#K(���dճ�qkru���8� �A�$��
9��^ 锺9Hq0JH�&$J^,�� �pb �BH��AJ6�F�m��Bb�d���]i		����Ɛ6c��0������ųR?=� �i�d�R @� CQ����.W:������1Ѿu�h��j����ն��!w����eF[z��	���xv�?Q�[�;џj��ܴ,l4��z۴�K��-�����������I���=�G�nn��ߑ�S��i�*�L�j$�yy����'��7�\��Y���n�r�V��d"���7��P�i餆p����՜��i�d9��Xд�����UEI*ۘ�x����J���s��˥���{O��ǟ�QRG��s��uf�μ��:WX�Tc��qq���qŔ�6K�˺�i���թ�v�M�g�7R,X��x�4+nYe�ǄTj�������]��7�hzMl��k��ŋikU^͗��l�K=e��u��WVYjGضdbh/zqS2�vKŪ2=��-zQ[�wG��J��${;x�Sk�jL�,>|ǳc��,7xY��|q���uu���z]�9����6B�AJ:��IK�������g:���Ϩ�U+D)�Ҧ
T��eaV����1SZ�+F\�-��4�.�.R�x�H�y%I5VP�jk((��j4E'4@�B$#G�O+I�ʸ�p�*G̳����y����y��H�(���Hvl1m~Mj����#A�`Э���L�ܑN$#Е{�