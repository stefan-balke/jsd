BZh91AY&SY��  V߀Px���������P^q; s���u������M0� �h  h �i1L@�  4    Jd�5S���mM�P�� ѐ�ɦsbh0�2d��`�i���!�*I&�L�&i�z#���A6������L$�R%���諜$���K�$�)uO}�U����%2@�A���#a.�ñ�yo��]+����\��7f�����7��!)R�(ݿ~-(�c_3�ܗg�=��\E�7�����!o[G#\�
��[wgj5N*�Y�DL����	��f�|�̴�c��]����
�R�q{��(���t����BX�����p��Q*��� �u[)j*��pCP~J��VG\��H�˩T��L<£
G��P�{��2�d/O8�
�!;ε���E�d�119ͬK�bJ�Ϊ�#X��H��ެO���#u�r�@�^��&]��}uZ�_5k0���f[c�p���I$�
 c<���b<}cNFLB��b��آT�ݶ��KEݬ�����1��Ć�Ȏ���H2�I! ��הs!
"�4���/��W��l�tZ��l��G��88SOΠ��G� �"TO ����3~]�H�`����������uܽh>�6�	�����f�P{֥�=w8�q%�qKCM���:$��>Je�I��1t)X}#e8�<��qώE��70=����Zd�����qBʈ�;���Æ}(pQ=z���:sJ��:/*p[m.�n�tc�*�|z�4���$�k`��dc�Wx�W&~���ɲb�.�z����f�EE��u�|se��Yz��r�Y�����m�N�Fa�^���px��q�?6m�4�7�����Mƅl�{w�EF���M���ǤTt1�+��ہ��95�/�L�5�5P������}�־DF���y�HXb�����D`g.ƛ��f[/�Tdz��k�k���lwy"V�w[��SSը�)7w�{u7�K�]�m��K��u��u<�S%�W8�%GIJ:<�a��K�Ms;&gx�hHӯ��(V�G$B"��Dn���me�%��^��$08�$��xsYhLG9�l��PtQ�2He���av�L!F��w{%ݕ#W�rjqԕjΞ��=�\ɺp1�7�����U>��~�֨mQQ3�3a���"�(HHW� 