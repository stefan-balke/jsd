BZh91AY&SY.�,w �߀Px����������P��v�9\4і���B��OS�$�4�i�4 @P�L�  h  D"MDؐڍ=A�4  �40`��`ѐ��&��D�К�)�h	=2�@�<��hI�@�$�Q$�������L �B��
A���Y��\��b4�XIGsRr�@�>��6�<4��:d��n&*�����_=Q��s�2�*p�aw0	&�,m�Z�a�� �b�����:2Qq�g^2�A�=C�ķɐZc;ƶ��\3ƒI+ki9�J��G80~h5�d�9Н�0���ۜ�ku3[bYd�f ΡB�4x�3>��e���K�A7(T�n̛5�7�
U>�b$��Az�n�I\���h��-W�����ʄ"�%1[Lw&oU)h,]�"@4�JZNr���m gCS���,*
�����ט��cO�i��1hu�K�f�++a�I�T�����,V[+�v�+aԫچ��\����%���rF˙���k��F�dj�Yz՚
Tyu�I�RɆ�s�61���m���j�r.}�;�JJ�עj(�.oan�0�V��4��ǃ,��8�t;�V!�2�2�H�2��`1�VI$$CZ�3�����*�j|26����_(�����%����N���n���C�����$	v�I�=��#�CNn^S�LKS-�94���4�'�C�Ё4��*Ƙ��5T�E=A�	�3�|�<5
�� ���C3ܒ�B�C=�/�Y��Q.�����|mD����;��dy��O��۲�m��j;5haA�!C��pj��D���������k��gf���f�u�5���61�Jڂ�g�~�4��vbȴ�LP;�'�{���)���r��9��)��M�
m!A�H�K���d	XL�KG���rk2�������� ��~y��l�m���i!b���$ ΀/o�z�h�S�}�P�.:C�oH���&4)��/��=�RA�� $�p(!D�P�!�{�E����auJ�XR�p��l�ѷ�~�'�Q\�]g:
 �I�
�r[h��4��7s0���%�w�3���9���'��M�3����(
g�*�Y�k."��� X6�3����q�B&=� ��l�^AY�����g,E#�3�H	F\f��66P)5�Ȱ7Ժ�I��St��2V a�N2��T��F^��[I�{�7t��X)5����n��ݡ��mT�m�mH���0hR���rE8P�.�,w