BZh91AY&SYmÛ� �_�Px���������P�s�-�84�T��O�<Ц�4ɈdL��!��hLQ�@    ��SS�M?S@@�� i�4�4�A�ɓ&F�L�LD�CSi3H	��OS�y@ ���yL	�<�"AD��A����#J>P��
I�LI�@�M��ċƅd�0j�R7 ]��p�i3��h�ZQ}��_~Q#���T2��0Z1
gE�%<Of���l��F5'g)��Ys-Q�j�a�`:��41U/�"�!*֌�	 �zN5�7�����Ly}����"�p�G��sn��eSRҙ���Rb|��Eq�d_
(JH���p�{g'��U�I�(О25"AIKD+�UJ��Q�Q^_��FT�h���r�V#�>�����m��@��z޹"J��M!	K2I$�Pg?!��,�tp9d�������n��B5�
��IJ�]�.�!�l��D����YKI! ���፴		BDfי�_�[Յ�/�c�l��j�	�e�(,�����&�GϷ�\RP�o�F!􌗕K�a���(���X�`��P��V��1��� ��0:��wi�S��k����z�2٤�{j� =Q��3�@�TPC�zY�C2(^�A�nē�@�kk�kw0�uqj��.��TP9\��&s�J��+��z�C����5+�`���%L��^������q���(K�����8�YA%�I*��z���o<J6��ж�~���֦`L��0��L��˜H�P)���(
D�3"cc�)�hԵ�#*��i���W�}m�THc��,�F�a��s8����Y4�� 0�N�2	
l�665�~b�K����ap�2��d@F��ބ��>c��f��ԂC�&x�>��3H@��m7.�g\���Be9��0�$�@��a�׸Ba3�yc��.��wECHPm9�g�p�6�љa�x��*�+�g�Y��X�BjN�
SD����J�B�����Z����
�A�;���F�g�Q��b� ��l��-Q�����6�&�K]�3��`Ю��m�.�p� ۇ7�