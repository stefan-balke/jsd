BZh91AY&SY���� �_�Px���������P�]�&�����T�&ʞP��橚F5=@ ��(Q�ML�P 4     �Ȋ�SShS�0A�S@��M0���a2dɑ��4�# C �@Dɔ�I�Sj�M56)�P  zjz�R�g1'�!�   ~_/��# = ��
#H�E�0��ۀyI$hJ��ar1�Q�9T4�ؖ�M�QƏAּ{�G�w�`ϝ�0Z��̈F�QS���lu.��s�9R��_q�䡁	�@�&�X��k}(���n�	�=	�I��~-5��X7� B����..#T�������Qc�S����p�'�:�b���"#�DJ-(����BK\���S���\#���)��6�;,�
=�BaF�Z�G'u��P-��#T9��tأD�ڴb�0ЭW��	HBX$�J@�qC�1�r�g�ˑ�J�#����ThB�%m&�BTA�D��a���&!a���A�j�P�-����e>��ᣳQw(L=>^��
�
)GU߅EA�����4�B�!��𝎠Rz�}"��"GP��Zf�0��K+1��|�!�
���VlV6�}��Hw ��佯���ڒ��(/����
	�X�Im �d×�� {�ƈ�c��d�E��ƍ��#��9F��9��&����D��� �Hx��.C��>���ob !��$��
�=�� y��d�N�R��#�<��g�R`�{�d1�P:Ǝ�#�w�����6U�ж>ݙ�Y��b�x�:�{ana����i2Am�[D����<iJv��";֖$j�h9v�8�ca�a���p,	-�Q�BA��R9��*ةyJ20I�f�V�����>���� �G�A�*��@�B��;���ڄ���5��7��� ��{G�C��̼ ����G�9��Ϗ��*DC� ����~H1	�U�N'Q`p�4�1�䁜��2#��Q!�e¿l7�=�EH"����ĩ*�]�7�ACDS ���p�m&�[l"�É8�1q#D_r�m#g�M&.B���
@��B�vk0X��c���G��Ը�d�API�d���ܑN$.�)=@