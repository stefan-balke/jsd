BZh91AY&SY���� �_�Px����������`_<���A�@h$	Q&������ �   	@�dFS�mL� �2a44��& �4d40	�10��5Q�h4<����=@ h ��b�LFCC �#I�щ���L��M&�= � SLjha�hI"c$L�"�W�����!C*�uI���?�*�ǆ	#8Ю2� �F֪����ﵰս���j�z����ifYۆ[!W���3"so��]JuRi_ 
:���yw�%�����gu!����U����|`�K �)���"�q~�ZQ�!����GށȜ����q�A,0�9��Q�1ɞGws��fX��=Wr�D< %	�mZO���:�&��ꆅ/QQ��߾+.l�5*�,����ěTe��jv�nX�*]c2��f�a���C.���iiXt2�3��w�2���AaR��f�NX-�d.�%*a���dˬ
d�Lg50��M^�D�Y	��wb��)"�(��RG�ȣe�y_�¹�L��3�sl�b��\�ˤ[��b\���P�[Q3zV��0�f��Ŕ-$�Noۋ7��:m�aEك���;���)Lk��Ϩlcc��m�4m���<4.N"9P����*Q%�aH��*��P�w���E*�P�,6#rF�Q���;����=��lh��aشv ���&�&s����7fǐ�}9q���ġ&��:8�b��7��SS����<1 dj��)�W__���ͅH�xT"!��ӫ�<���R�I�]т�>��wl���{N�3�(�hX�h|��rh�L▇Ǻx���S���$�v$�#��k��������4JZ�\��g��Y���V�K�~L����c��B�ZY���b��5LB�ȷ�Z�I��a�U�73�pg�a��8=-QDU�1yv��U�J���[;&ƹ�03/�z����^�>��Z�ǔuy���w�Y�(���D�]�>-�)�c:^�.r�^:���~,��ir���n�,X���m�­Ye�n�X��u92���p��e֮ʽ���.��,�7�e,:��`�ej�ua{p��F������"�,�@�3��iD$2Jt
X�0�Tdz� ���u$���k��̓N7��u#��������Xs����w$ܚ^��9�t:��e�W�i
���qvn� ŋ�p3��n�:q8LR�aNne.�#�]X/M�qon��~��Jd+`�Љ��nY����HF�`�7M�aQ�:	�/8.� �c}F�vP��v����T�>5˥���;�y�[
B�ͳ���o�]s���U<�9�~�ԨlQQ88�����ܑN$>�x@