BZh91AY&SY!xm� Q߀Px����������P~wcXa��h �EG�ڦ�L�4�bd�L�1 ��jzi" �     S"�T��	�d���cD7� ba i���&L��L �0L�0�D�d�bi�	=j4 ��i1�:	��@�*.�@��?A�җ�U�Hi@2M��6��i%xЬ"��ТT� Y�ȼ�S6]]�[�ef/�^M���.+e!B{d���r�� �"6�$��Ի,��[U�X���=܁ㅵL��5�u�/ �<�z�fz����j4V}h3[Ns@�Z�NhP�f�x������H�{��0c݇��(7����#^��������&'m~�J��v/P�*w[F4w�@�ù�sL��@�ZEȳ�*"V�)JL�QR�(�U L�B���3�J�ZSy�Ae{,�w�eyT$���$�ql�I%��"�F���6���W��THG0��A���%����`1>����r��xM�N���bB��I$�D�G�@nI�r�s�ˑ����0�!�A�G�]-&�B)��g��+���"�$eZd$5�F��6��xF2o���W�.�Xt�=%��1O(
|�>Y�F���:8&��C.��G�Q�n ���gǄD(�o�WZ�
�aB���7d!3����!��C/
�l 00+Ns<�H� ���`��^#6�IuKڀ��6n<hI�06.�+!2�g�C��d|K��O*�[�Σ�Ƴӆ�����˃TP����!����"��BugY>�s]�xz̖�BCHq��.�W�}�d}����LP%�{C���s�@4��Ck5�$�K#�����y"(m�1�����EiS]��03����ȶ����ж4@8ʼ��#�Z�.-��@�Y����4�������~�(�Ib7��a�H�$]&P�J�4�	 0`0�>Xd1]i�DA��R/,�����$7I��PRh�v�H"l��~�׽	��W�q =G) �@`���VH�4���=�w���������A�hL�A�9�Ą��� cs�Ā�$L嚼��t0�/�X0�Tm: g���a��8�LzQ�p(3o"�"����bu	�;��@T�M��A�1�I��2*-~\0�n��,I� a����K��j�>-F-&-G�H��L/h7��Q���������5KZ�ٙ��`��c���rE8P�!xm�