BZh91AY&SY�UU� ߀Py���������P�Yۤ�7/nM��IHj�&�M�5?T2 =@ M�&�� 4�C� 4    BdFI�i��L����  F�EJj{Eh�4F��A���E B4h!�j�i'�j�h�z�H��A��0�TdE.C��$�DH�{���iI���d���3�͸���A��0��A��u"���Լ��t-}�#L�iE���Z�=QъH�_t�_+��7��7,�k$��1���z��^��4[�ȉtu����(Y�������Ht�� �"'��P薸�OB����R� ]k�(�.��Ҽ�el\��K����h]H�������dF(�]j٦ی��1�IA�,�Up�GAq�f�p���p/����NtՃ�*떕lY4h�tCi]*�5�9��C>�,�*O0G�U�``,��� �̈I,�BR�14��@5�D�]j勳�=g$h.:M�����p�UWغ�1�"��ZBe�
��jH���Y�b�����
$�*H���	�61�����������ʗ�Rn�����w)��QQ%��m�n���Rt\�K�d�.,ʈ�a#rFƛ(�q�ʨ�P��H�a2�[�lm�s�����6f��͆�\����X4��i��C=s��`���UOI��a)�;�Ȋk�y~un���;̭!陑�.0��̴$)��6{�������^�/�!C�D) �O4JZ'�^&��0�R��f�D���C5����ɭ8V؁ m@Z�Ԍ��������#ȹ�	���o�-^�t�-K;o	��#".+��Sxch�.H�{�L�H�4X�R��W�s&pߝ���^jp{�H�1'"�7�o9�)	�o��IA�T���W���͌
S�ӄ$]����-ş墸�R���`�hJCl������b���"w�Oeڈ$9A�H$��7�2�k<��` ]P�m�:���=
@��!<���h8�Z˂}X�u�^,�s�6�t�)���@! �o�(�Ab��	��I�U�W�IU�f2/"�I0���$�c��m��!D������R*������#�ֲ�����fp=+�|��� A^ô���#����X!x��P�(�A���o/^�o���,D1T!��A2�%��&<�`�,A��<F�Im��u�2⍂��%T,d�q�DEq���d�ҡ�n�y4���+7,I���]������\�����
x2z���z�505��Ix��#�����!=�i[��A����+@rcw�]��BCQUWx