BZh91AY&SYQ��� _�Px���������P:k.�〠 �4��Ƒ6��ڀz��@ j�!j        �������=H�h�i�	�&��0L@0	�h�h`ba"@���S�hI��24h4 4�L�Sh�! TH$�?��9@��
�)
`�&�����x�Ua`h�jNQ	��ۙ�f��YG���>S�Z�RQ?m���tb�&�M"�����b;��3o��H�]k�Te��G=Q���A3~�S�f3�x�kk�� V�7҂`�&p���2.OX)�!���
+����bI#���a¤g[:*�:C�Nk�*\����o��(�p�^21��.ʐ�C�(i��1��6"��ِ�Ɍ-0�@�"��R-	8�������C�%���h����1��)kh0Q�+bR�1������@�a�/X���uaF/��D]
���I��<ޠ�TF��,�!Eh�"S�iBV�!
`�!đ(�M��##)ykQ�,ڐƢK1���	cF�x��c&�z���<_�a}]Q��7L�:pY�0|�&uo�=A��a��D�-��ФJB�]r��b�k�N��0�F ���\���r$x�@`P�k�U.�P>�d � =���eԾ-�%��P>�_$b΃�@����мl�4�C2(_{ ��[�I�J��ٕ1�Ym�Gt(:�.�#��	��3��A�"`ֈ�aJ�#��U�x����l!�%9�������aq���(K��g�LqL.�D��I5Go]}v\	�T��h�腓��qE�5&��1��Om�7�霬�'G�#�ɓ���V���z5-mʼz�� 4r+���ʁ��u�%�*05�5BS��+��5�HX�[�L�ұ2 �!��;�vH�`��̂��eI�*��U%FJ5g�|�(Ou?�p.㒠q�ӊD�#�_e���p5�����B�xu�6�	��<��$'���a��!"bg�yc�s.�]�P�Nhǈ�iQ�$8Ж�2�2ݞ�V]�����,N�5'~����h�8"�Ҵ�P+o*Ծ�Xb�)-[	*�a�'�^�/���߉�I�� ��2؎�H�дK"�{s���pT�˿vb4�N�����"�(H(�z�