BZh91AY&SYO��� �_�Px���������P�w\�Pc�#M�	$���h�� �  d4h4J~�T�d4�@`@   BA� �����A�i�#@ ��b�LFCC �#I B4�1 �z6��!��4�L�r/D�	�!�#$�)�+���U�a�1��)%����=��U���4�#2�!���:$f@���G���_O/S��-N���_�j�N��'����,�P��D§'Lm�&0J�\�y�Z�����>�@t��03&�c>�Q8�ԑ^��}dq%tP*��-��x!)g�h�H�(��bbY��3�K���!F�4��~���^؍Vڋ�]����頳�*2�9H���I"�B�+!�"}@��5e�[*�i���ɜV���i��A�z���h�i�ɻ�b�)�	&mM�B�X�W�+P�Z-���K�l@�h�gX�l�h�РC�'��Ê;B0cvu�5$H�:�Н�MG�˦��+�žt��,l��Z��5�l���҅��Nq���o�m��ĈC��:>0��.ޢ9P��璉R�-vF��K̟���ڙ.S(mZF䍪c`ۊ�)#��da��kE��
�d��L�+������r��K$&ݰ��'�>~�Ws-���n�:���S�Y���J�������������d�����ㄎ���f����+{ѣ�Q�hX�9�s���r�LG0��U�d��Y�$�IbD~��ƄV���|p0Jo��;��|Z�����Y�e�$�.�gK���s7���dE���s�t�q	��(x�X�_VO��8�e;�MsOdTJ�l�F=���Fet��hg/K.�����TG~�j�غ:���9�n��1m�;����&����a:H'��� ��ᩀ(�Kut���V0�_��R��x�芎Y��lǦ#���=��Up5:���.�&*��5�_s���ۖ�8��ts("���,HK-C�v��F&��M�4*�د�Tby����Q[����%n��n����,��̗);���6�1a��g���[�^3�Q)�[��2\�^k����=�/��|�NǑ��'���U+T)�ԥ�T0�Eʶ-C���)�����я!�Tq<�%�T�ۜ��j�;��7�:^�GV-Zt�4hT�C��.c
6E�k�q���~nJ���Y��m4��%̛��#;���,{�rUO�|�-�3T6���y]�0�]��BA>#+