BZh91AY&SYt�+� _�Px���������P��p�!��4 	D&�D4�G�f�@�  A�h
M��      ��F��RmA�?Iꞡ��� z@`LM&L�LM2100I&�&�a 40�Mk�%q�%�H�	�B�W�����/� �B��,!2��E�n��)�a4v�T�Y�7|�z�>^|}�c��kZ�;ar-K��B!M5F����`�nzR��@�Ύ����6�WS�+�8)1+/ܠc���D��a Ą�mzZ�H�][�rau�ȘN�ώו�-m�n@�V��	34��ѡ�x�P��m������oyp�!4��Z�'0�������]ԴU��.��k.�qT����o�*Z7���g'A��ۢ1eDy���I�N�#X3��H�Yhh�s0��:P),���b,�YB�:�C$���U�q�Sj������f�7K|�#:�1M�n��5�%x�4bՑmp2I+����yܽTd����*�6�d�R����(��@�A%pLU��P�AR�6�Et�RFQA`��*RF$i5P�A8�^��plcc�m��B�>/|������#�
Bw��^�$��q�Ã=wś�+$0TD ڼ���Q66���UzoEֽ���(���αj���f��eކ偗08<kgO����%�8aJ��7t��D*�E��c����:�a�&]ܻ��
��g��D�#!Ԉ�����Q&���'�uw8��߼���<�4v)�-�o&��]|�s�R���Mq9��S����I>~y6�J�؉�Zt5�b���>XL�����d!�3ڒ~�cۊ�{D/����Z�K".W=N���˥��=�Іr`kR����J�Y��B�c'�o��u*
���N�cA��^Q�]x���cG��=���(�N�v��c��<���^�,��FX^'=v����&�v��e5}6���Q���LP�$�#�˓F�D[��Ե�Ӓ��6|Q==�Q�e�W��ቩ��7�[b��se$�܆V����_�`"���#���萌K�#c#I��Ҧj��/��#α%�KX�����tD�lyQ=���E7<�ې�����A���n���gc��⥡�ou�qWa�Q:�h�k���+�9$TV��6yz7��w�|��������Ӱ�U+S��L�ʷVuM�6�[�����v�V���u#s�x3_"�
ӫ��&MXJX��6ͦ�K&�ŧ��6���樞8z����p�r�0���ӹ�RT�س���4�8D�����&�"�=V>q�U>.������٭eN�n��w$S�	N���