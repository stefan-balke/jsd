BZh91AY&SY�@�4 -_�Py���������P^�s"q��vP�A&M)��Si�i��ɱ@h�&��Ji�� ɉ��0F�`��55MS��=L�Pd�4�ɦ�8ɓ&# &L �# C T���5<E=�=���b L!�4�IS�"Ȍd=�Ղ�+���*�q�.x%��T4� �0��0�Ö�CI\e�F����i��������zz�^S�P�yX���Z?QY�ƅSUPD���0ɡ9ə��Vl1sh�<e]02&2*�W�q�̦e���R��Q��l�J̧6a��0�6cd���sġ�|;'���@��x��FH��9�[Lv��wmJő˝DM�\��m0��K�h��3C���P|�螺 �ZD�g Y��^d=�Ζ���Cñ�VU�����J���t�g�ʤ�!��S;�$;���u���"`�E�E�Vf>��zC|lc{��I��5�<�����A¡@�&�%B�0��^]���LJ���j@��rF�P���2�UcE"��a�lm�0�]1�{�/���mOqj��ӨL����z�}�?_e����6\�����:n)<)�3Z��3�wuP�e����Z�0��I����+�W�W��q�\f�z��,k4;k�s�s��$���I���&.��J�x����l����0E7Q6�}�)Q(�:�=Բ�k'��T��Fud5>�������.9���N2��AgT��3��K�[Χ^:$�)�v2j��,X�U�8�21�+Wp�C_V�ഩL"'�g�_���i��1�ik6�;e����b��7����ͬ�дd�RW��*� },�r��f�T�?A����ڋ-�xm4+ŋ_6��J�T�H�Yo�)��"����O-Q����6ke.�10)�'"1-G3Bp�Y� p=c��*xc,HHA���!`�Z�w
fV�/�*2;�ȵ���i���$�ӵ��yX����r��Ӓ}mm�KR\N�:������r��B��Ǔ��d��#\��JRi����������̟3r�4�
�W¦�R�){\�����o1S��~��h�9��S~W2^ľ]\��0�-�M8��k��J����h̺2�G$^[1��↶B��ͯ��d�S8S�:H&z'Is'I��x�If�=|4U׌�,ަ$XLzF���*�-Yc�rE8P��@�4