BZh91AY&SYG�0 k_�Py����������Px��GX��@T%I2=F&��@      И)�� 4      $D�H���?D�OH�z��d m�d2i�# `F&��4� �TDh�F ����CMG�P�Ѧ&��C�@(I%T�]!@��q��M��Y�H�T d����p/
	,F�q�ah�2���"����:8g�ӥS��w}L�!���$�7�U���/L@��R����mfу��mSo���ớ
rMJ�X�d�ŮM�̮���wT�U|�3\�c�D�+ქЄX��(�R�0f��|�{<���w��@4��])������+o�|S�w������IwB�E���ϼ�wY�=��;�P�dҫݳ"uQ����ȵ0�3��%��ʀ�)�ܬ�su.������j���&a�&�Q2.@�t9�6r��i�*��蠢���1�@����j��e"�<�rp�C�߼�8�lcz6�n�=_�wUGb�enUp�S�k���*K�R��KRTxv)5���D-̐CH�F�`1�ALd��avjg��cCa��cT����w_<�܇��
�+ǪFmj1
�9)��Ԑ�+���f�����ܯ���Ƀ��c8v�x,�c
퐡��˷�;|O�<OD��E ����n<�h����U�MG�>Y�Έ���|D|{Qh���8���䑶=�E�(J�ּ��d�%�RN�������fݣ�Pr�:���TT[��4!��!�YEm
ll'�΋�C���5�G���c�iS��o;�i'�&É�Sފ�W��~����$9�5�J�p�:z-�c�����	���6�i䗈Ht|PeQ��B��H�1�]��\�#t�B�:#�̞+Z�.�m�i�S��s�������5���+����\\!\`X�kh)C@�7L�1�D�Ȁ $�h�D�m� ���"�Bl�X&�]
L,z�AK�J�5Cպ:���,.����P�k�����ڱA���V��r6�O=��6&%��g`eS�irRh����Td`�u17#�&bo�\8%T�_�����3���kۿB-H[!�,4��UX&��Yɗ��-b�%��3���r�}�2b�����J�,f��|�#?��74��3��F�Vq�h4Vn�ȩ��Y��9�o����i<���¸2���H�
�Y 