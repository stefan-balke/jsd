BZh91AY&SY�3u� _�Px���������P��h�0�%5 �)�7�A��M43P 9�14L�2da0M4����$"5!1i�G��@�!�S#`LM&L�LM2100	L�&�SF ��OH ���S��I�i	D$� ��OW�ts=�Z	�,Be5����o��F�B�&V���Ԝ� B�@Z���9r��>=r4r�����]�� ��ɒ#���r|��vڅ0��6٫T3&��N^m��7in�����ui^A�z�&j"�p��Y<������@~7�@�C@��vF/d߯���G���DA�a� B��b�ĭ4�>��\��RLU�E��C6[ēt��m쬚1Q�L����?$�!9a�q�5͌D����3������[�E2�ra�7P���	�4Xb�ELj���M�*=�!�SW��VhOU�j�p�e�er3�K}ho�74m�{6�|mMMq7\Q��U��o�����"EQ.��*d�ע�&��Xa5*�q:��s���wAmu��s��lcx��m!A�����Itx�B��'�D�D�f%P8Ș�4P��'U�*)���#k%�������$s�#.�oB��A@�&�N� d&fHi���K�3��BKV��&P�&<���M]c�s������Ħ�`
Մ��"���J����5IC
�t��[s��l��F��f0G��m^p�u��3IH�i��^v�]��Px�!2�^��l�ѕ�$�;@G�B�Ffpm>T
	�0+^u�I�d3a0�����a*R�2
&5cB�uݛuc!%�tojhL�[�GBhC8��&�
Typ �^p3Ϥ��]�(�3&.�����~@j��F�L��B^���z�L��A���$�GgU<B͛ʈ �Z)Tж�n�	�%Q���z��@��Y�<M��[X�`�6��Δ��~�h�d�A���_����N��6&A�"�[���Ȩ1bUTf���T�"��Pw�PY��$$#�Ia���e����h���%-�_��|��Od��]�8���8�$1��=��� ����/h�;�>��hL����HO�A4q0�AǻA0�D�L�Ņ�ahq�4�ciԁ���$1�7�����ٻ~�"�������P*]�Qu�*��2f��`59�&���H,�h]D�)�a� �/%-m#/W�F�Iyr�6��R+6��	j� ���Ղt�Y}��&�R&�-rE�.�p�!�f�