BZh91AY&SY�^X $_�Px���������P8^hC֔� J3@52d��h0�42 ѡ�0&&�	�&L�&	�����jz���z2i I� A�����&L�20�&�db``$!��h��ښ<�� =�e,�yБt��$Aۻ�:�6#�dhT
��M~C�f��� �A���Q#H0�1|ڎ]�t�Y�v|��`�T�'Oc����2-�_0�*�8��v�Vn}�p�X��R�<�"$(��N���A���R4בДwҵ��f�1�2bP��qA� nQ� �O�z��L�����1[��Mt��Z��ȶ߅R�e:�
ٲ]�2�-�x��zc�'�$L��;J�-J�W��g)^�+i�+36W,pp�X5�`]�p�TEM�b�We�$�l&�ۓ-� �&�� ,�H�wB 4v��z<]��9�61����m�4(C��4w��Is�#�
��Q*Q%��v�6�y+%Gej��L`�nm#��2����4PP0�s,��Bm^際������G��QA��!'�=Q��a�%�^�ڃ7}�f��z�g�=�p�$�:ɱcUuJ����.�P@2	���I{8~6�ƉA5 0<&7�y�-��@�$Qul Y�z��U�#-�%�L���捌�>T
	��7/+!QͥCǹ�A�-ڒzh�mzjm�b�u㭻E�".V�����ˋ�1q�(h`kIN���N�/t[J�ı�a�P���mI	ma;��<�2�D�)�.d9��i�Z`�q�r]���:�k�/�y�x&r��й_���������P3/MX�"���X	�Z�D``i����Z\�dپ��P�T���x��:
�������5�\� ��̘jiNe°�ٜ�5HY�<*��|�Ą�i{It��!Y�2ÜʓD4T=�D�l��ݙ߽	��]�10���iH��zK����r����#����y��6	��u�d�rhY���&��cg��
�Ĩ�y�X�:Ϙ�:�4\���AQ�聜x���MR$��2F�h�*3w|�XEq|M'=�X�BjOx�SpM@d57�U�rAk\�%��%*�����;�F�G�Q��`}�=f����)9&�J�����my�-ݙ�уB�A�ޟ���)�
�j�