BZh91AY&SY��� _�Px���������P8o1l9�� �UO(`���       �MI�'���i�� �20�L�`�BB=G�4���  z `LM&L�LM2100	"L��
O���2e4��z��SQ`�� � 2 ������c��E��He5�/śp�dA�d��4w��R1R�����k���ى�ν�_Jen����<-b�[�Lm�����ꑊ�ʴW	��(�Q]�F �����#�\�4�@�r��n��$R�u�B@�p�}�PP�d�T�����H9$2`a�e���Ek�X�����	k��,��m��\��0�������\]1j�L��Z����T�r��W�D]�'�8�gZ��j�Ū]�+$��_2�"5@��F��uM�th�
9��vw���B��RfaUV,�bU?�61����m��
��8��Ix{r�Hw�tJ�H^�E1�`mZF�j���S�y9a�rF�L\L�ʨQb�
���ш�a�g,�M�}3˞<fl����P�$�g��pe$���ȂZ�q�6xmJ4�����!4��ܱxC�I�	�BYu1�{�-QN����"BȨ��2 D�^�{}�v���/;Q��})�K���w$u:�E�d}b�Xe��ԅ$;�sħBI��!9ҪM���i�s&!ƹ���ˣ��o��6�5Η�U�yÍHg��(\��q!��F�B�>ct��myE�"��s��>��?���02G�� ��l�ˌ��VZ�6Q��H[�,�-��D�"p,�Ӵ5}J���`.\�a88>�1�������a�D2/X88e7$xu�28��6�`�Aa�/��c��\L�nZ������Pd\��)rBB1{	t���XgP̆`�s"ȍq1'����2��D&�x�}���b��x���#�=��X{��㬸 +�v�������d&)��p
�P�@��/�'�겇3��-�b�c�c2h c��1&t@l�jEپ�2�V�M�;K�)�fZ{-�M"�[��r�5�WZ�hP7в�(2=D�[�I�p���.�H��gq��aPmg�D�hD,`1D
�I��!��p�̵���*U�1yP�2i��T�rE8P����