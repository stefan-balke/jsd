BZh91AY&SYS_�, �_�Px����������P�rf�n P (�LBM���i�4z�=	�@ �@�h�        Jz����L�@z�I��h=@  �4`�1 �&	�!��L���&	O50I����Pdh �Kɡ'�P�D�,H?�9	|aZ�4�`&I��|�1 �j#$00l�	�V12�\'c^�C^�N�S�&�e�8]n��	��J'���jMYFn�a�Kc9�둯+���'X`R>7L�x��t�넊�i���Q"��#�gE3&礌�>�(��{Q5֍@DpD�����*�=2͋�D�aω�QUQE��y0��+(G\�Mv�y��~�n^b�M��Y�G����-�꼱�ae�Q}$LO:_f������d�fA����)��9ɸb�V#pL1� Z��P
X���f�<����n]�H��B��R���i�JK�*5A3��*(�E	�m'C��֒�`2Hr�[�PA�I@�٩XK�U4���h+$sS�P�b`ޠ@�Q\�E���&���-�XQE�*�I�c�`u荻	f�����D��3k�I�)E��ĢQb�����+�V`Q��-"�!#���(�A;��@���ETI�Ҭb��I�����dNaaP���S<����_\�Z����YL(H��<)�Q���ʱz�1d `a�/�ѼTE2�����f`�G��V��� ���Gy�ۆ�P4B�^X��:��e�%�TK�|�����B�3s��&4ؙ�H��>�S ����$�J���f4�^c��{v5�B"�V�qj��@\XqMd��0k��U����̃��Q�D�A��f����H���X<�.@)�j�$
��H��-���5 �^=�dפ�9X�WM~���y�(H,CF�1��u
�ኚ����Z0��[�^&���[Z�|��^?5k\�s!��!6nz;�9�[��� İ��A��0��NfaXnyN�0&��� $r�@��-��Dп"�$P5�Ø��5:��*I`�d@F6���	��Q����H����v&Ղ G?|���>��4&v�� ����&�@��� Y��L��,:N����EB��i�8p$@3@]�-q��F{��A�nᐫ����#��, D��$���Ġ
��Ah``@��� [u�����Kd�T�����#/'͑�I�q=d�&���h
E��e�P�� f�$����ʖYo��ƃh��j���rE8P�S_�,