BZh91AY&SYs� _�Px���������P����]B�� �EO�FJzO
&#@=OP�C@��M5)	��L #CC ` 	�M5��@�P ���9�14L�2da0M4����$H4��h#ji<�� 4i���X ������h$@������2Щ0HL��A���+@�CB�e�@�9�)�@�h���8�q�ǗU���o�F�Oi֪U4R�*B���������Ԃ�dö6�],���Ӽ��D���6�;��ێ�c1�s�_����KI��+0%�9um�FK��1 ��sBB��	����b�R#���O��"����p�ֱ	�	Э���|�9D]gY����⥓�W�;��1:�%f�r�+��'�	VP�e4h����1�����F�l̄D�m-p���s�4X8D@F��`�lnJY�[�+b�����Ɉ�
E��{& 5�)
Y���"��Ba�8.o���"�B��)&��K+�a�#*�BK�lA1GA�ů��Y��q�����l��^%���5 �A��m�0J�w��pR[w����D�D���tK��|p�4(�#ZHܑ��J�mF�tB4�`�l��TT(^�((F�&��bm ص�X�W���K%���)7�����9���B/���/R4�T(�F}�����\ܹ�z�k�[����Ŋ�)�	}���g�z������.�i�A�^w?i��B�{A��	�^���ҿќ˷�������H^h���ʁA3{r��Y	�ͥ���A���I<(�mvUhe��՟Kv��B(K�<qj�C�Ԙ$�B&g�V�G�:�z����7�i'8�y��A�Ͱ4�2T�����>��d�4�� �IwG
��ʿ@]����������qE�0S9% ��1� ��]�V&ԅ�vkf�<�4U�^|7���+�!ys< h�+�{a����b\O����������F����PY��$$#�"�FPVY���̖�ѐ�2��� "����	릤��8
`3��JC�/+ׁ��O��q��F'|�5	��;b@��(:��4w�HY�L��iYˎø�B��P�(6��3�����Hs%�����\3f�ha�7��}�X�BjO6~L� � �hZ�A��o�vk��4e%��IU	),���i�=؛ZM#ȃ�Y�306 �cb�TFRD�H>�m|N�K���!��0hY��S�rE8P�s�