BZh91AY&SY��� I߀px���������P��֜ �F�Q�my4�b 4���h �@�ڙ�        	�@���=OOT4�M=@s F	�0M`�L$P�&FSi�I='���OS�h d�p0� D���A��~c��H�DhT���I�פ��n�Б�дLфHh�ڪR0�ϧi��˧L~�E�����"��/B���Y�����`4t|�H���Cn�G���xm�Շ��5ꑥ:îp���0��W���0�+�g�Bq�~�M�C+�zB/X;��@P��I$)�9�����ru�Fۨg���Wy��M0Qo�ϴ�bP��&�3\�ǐ�����.��q�h��A]wh<���K�ݫg���,�.n�i" 90�j����Y(�&	ra���kV���x�Z�10�(��s�D�cJ0����ʋaL�z��^� ���W,�i�j�,�D$�&��Æ	'(�B�&+dc+l6������`�B!�$�PT��X{D��D"� �l��]\,��*���� \{D!�@��p��Q�ǦY�����p��������7Ŷ�h`!�|'��>zK���T)!�|�J�Iux����(mK�Q˪�u��
���n=[U�"5	 ���c.�m@B�����k·�DTDD���Ut���!����w�)2�D�?���ZX8q3j������Y!�H��n���$�y�b���b��U�s��B�X�����K�j#� `n߷�������
�Ѥ��A �-;����b�x� �T@�/[R0��4��IzsJ�6�I/Dt3a��	�01\�D66&A���� @���z��t���CepH����ZV���*#�l:Z�!�%��d�Bg`���S1VI�����83��hq[x�$�b��q3وV�����i�`h5�� ����z��$�D2"��F����~^��yQ!�q�/�;J�йH�$oY뫪���'0""d�t�AL�j�D!Z�hԮ`���Ԓ��< h�'�}�� �℉f"c���JG@N��FF��J���HHF�&0e����h��-�ߕ�xmBxXOZIv���T{� Db9���Q�� ��a��"��!���2{���r�o4��$�	$J��^���@o}s��䁛���T���	[�3&3s�)��3�Ft�B�����ɺ�BC���.|^��-��R�H�*���dT�0��)qiz��1i4/"WY�h`lH�Cb��+�s�|���3�2S�_^^A�f��E_���)�Η,X