BZh91AY&SY�H� p߀Px���������Py[z�a���	B&��L��SL��=M@  J�F�@z��     $$MQ��0�@   `LM&L�LM2100Q&)��ɀ�jz��d=  #G�׵�}T�$�Ii
'/�u�6���2hT�J�!Ms���Z �(*ʎUT��'\�i�݈���[D1����j���D��>�������{9��/Cn�_ǡ{	j}�K����8�r�9�#�n��Ȫ>�FRH��+-q&���*[�y�	$ZԄ\���#�oLaH�I�����;BbEj���2����\���8d���ԣ���ݯ�j`c'�4ί��b�ٓBn0�j;��	��AD0�4�\z!�-��%j��ib�Hf:3V��L:��3L2@W�=��TT�4b��Bnk��I�]��f6��
�R�A1�AɎ�\�"��և��Օ�ϊL�-&��4J��J���)L�ocm����{�v8��Iy8�B�w��%J$��Ci�Ӧ䍎��X�W+��̬�e�Ri�b�iAgE֮�`66�b�����L��/!�9ڸ�2����N��6s�1�Â��Pr��L|M�e��-=���)%z\\"�s�{L�8fZ^=Ʉ���Ǿ;�����y���Ԡ{JAC���O�����X�J���GM��>=&n��%�TDx�/��0�-�W,�q��?�ЪI�T��xz%E�o4DNV0���]���n�,�m�!f�)�b�V9ˮ%$3xE��R�EY�������ݓէv	14ֳ�i���?H�'�}��/Ȳ0.;)pu蒚QA@18``b�ɶ9`��8q�wrUF��al+�>����QW���Z>9u�,���۳&��Ӟ7L(STx�4�e�?�eDrN�܃��zDñ~��̛�hi5�30䋤t*e0V���3]u:�����t��X�$$#A�"�BƂ��\�5�����R�*P�����;��;�%D�z��gUD>5����odPwvz�oj[�{Mi�K���n30�=C(��a):������q����bv#��ɘ��.|��)V��i�#O
r]-��iE��9d�K�l��X�s��]�R����iLR��>,���*��;�a�~e~�H��{�N�I������M6����/�!G4=�qmr������x�tFM�w���"�(HR�� 