BZh91AY&SYZ��% r߀Px���������P�+�0��!#����5O�Pbhz@h   �sbh0�2d��`�i���!�HH ��M��554  �@sbh0�2d��`�i���!�*��$�(�3D �jz�ez� jnY}(I]$HP@�<!�lK�a�P4��MO��8�,$�A�a���R�H�f@���N��>�3��a�>׆�3�L�z�?{�gd�������%�c��+­$��Y��>�=�^�,`fJ8�lG�,z��(�#.�:�`ke��Q�(�V$RR�9n���)!#�q{2'e�����y�Jx8���u!�0Ft�R��ע���8��9��W��e�B�}�QX6-�Shģ��7B�3��3�jtJ����s�%y��ڇWj���*���6�l]lgJ��Fm,^�4��&M.]�ɉ�a���=���ܢ��5�,��cU�5�7�K^�v+^/�������7eb4k@���u�lc{��mz>���Iw�ʅ �=J�Izv)�c�6�t�l�a�t1�id��P�ƅ��E@ւ֊
�~8hM�sǊ�4s�<�q�K��_�,>�;x�O�X��ڵ�/8�u
��#PF�g�{�2����̌��D�6���H�����7����_Y���ć�R
�.����\h��=J+������LG޿��Եo�����G�|���֖�[�i�b�D�-�����TQ�0�"']�n�t����c��72�9�r�v�m\\:�v&�3�E����`�[;�����Ưe�0��K\���w'���W!���X���{����,�Ij����}����a��gt&��Fs��b��k�K�?�8n~�\I a|U$P,��H4���i���l&�S�Wh=��0�]֞ٓ;NI�+�܋�1Xk�,��]I�2���dD-�
;9TAb��$$#A���B�΁��`�#F�0 �d�7=�8��xn�O%��k��J�ό"�C����,[Z�ޏ�����iI�&Oa�a����/V�Dà��=�"�c~Q�{����F7������	o�*��f��"Ëd��&s�zw"1�t�C�4d�ʞ�u ��k&PsK�7�mZn�
�ޑҶ�dV+t+k����1}'n-�(x���fj��*���p.���i���	���E����$��I�j�,0���"�(H-}Œ�