BZh91AY&SY�v� �߀Py���������P��:A\Ud
p�)�i�F���      h	�R@  @   BA6�F�$z���24 4�2dɈ��	�����%4i�ҞLS�i��L�4 �zMK�J�	.�#	$e �
��?YА��hT&�X�jz����a �hY2�	���t�,����	ß�n���yf�hZө����t�Q=~����0��@U��^Z�ݯ[mc��U�=���9}��ݶ�\f�q�����v'a��0��f�,x%ޖ��r>'��$��߭�Y3T{��B������T�u��w۸�t��`�������f��[`R�\w6Ħ��^�R�bm���.���>��hN,nzLqixF�3��|qj�M�f�*�{��׎���j��6p�A"�M"� ��d"=��! L9�!��!�DP�*�5A� Sĸ$	�����Mju�%����U���q�����3�V�j0���&#&#4Wr���%��������T1�DW��i��b��.c�xF�61��m���B7�_�<����#�
�;(�(��w�I�dS�k�(�����3e6�F��u�X�Сl�PP0�n�\�@Ɠk{Oپ��}ͦ|���w��;�� �o�äw�	ES.J��a���vAN0IsO_�v]���N��2�*���9Nz= �s+���>�.�������Y��su(O���Z�6�ڟ��������D���q�eݩ�G�'tl�K���)L��2Bdgx�0_k!
3ؒ|.�gM�m=M���vU.m�т�Zn�SSƎR�&t�5�_R�E�g����oI��װ���D��`r�dc�W�k+6����^�-��w�y�(O��N����ux���6�^��n�*1���ϻ{	��/z׹c�O�{u���C�4�` BA �#����Z��Q�5�Cn<�v�AQ�c֮ʣn	��g���F*ם��1�U��k�����@��Ƞ�wı!!��H�j��>a��2Y�!���..�߱="V�6������)z�=�����Ap����=	Y��\��S��f��4�kxd����74�wzs2yV�ƚ15*���9rR�T�p]h�]�s�W�2S��-i�я9�Jf啙/ľZ���	�M��u65MCx�A�0k�A��Qz��e�Rݵ#_Ʒ�tԔ�ڹ��6��7̛���13�\�����ET�8L2��S5Cj��������)�{��