BZh91AY&SY��7w &_�Px���������P>r]lÎ
� �(�<4&Q��x��� h  ��F�  Ѧ� `A)�$j	4h=G�M1�h 0&&�	�&L�&	����L����)�jh�1�  �����)�$B@��I ~>��r�6��*Ф��2M| �M��1PЬ2�L0p�TJL�3!��Y����u����S^��jJ'��ǄjMX�ݹ"��"5�0�0yR}���i�2�,\b9�F^��e�5�H���w�lz�&�u�1�l.G��Y�h�XL=_��r�A ����d��,���3��wie�1=�j��� �g=�`Z�6䈲.�7c��$�GP�F:iY�F�CS�upL�
d^��..�����$�"5cTT�B�#b�*1,�1�MD΀Ø�V!18u"�������i�H`�C������n�"��UU��$���5p��6k%���p�-SD�L0%9�a�%��b�"�ʕ2#R��BZ�3�Il�PP!,di{)0�hy�M/�;0l�a�;i/�	Y��T�`0a5Y;�������������{�
���p�檮W�B�.xxb	� �]�n��f���b�j 0&	���p�)��*T�5��@����b*�_�����U#�捬��PL��޾B�!�����A�[�$�J���2N�-�^��Pnd"��_��At�%�"`��LKIN�w�����χ"�KWj�6�������0+���DP����ָ��7�����:j��U�L��w�$\��JhJ��r���02�M0��6�%+���J5�=�U�{�oI��@�W�q�����}����23̸��03&4�2�7<�(ȚB�� $qؠD�d���A/Ȋ$P5���,;�P�DCE��,%d@E�潜�Ou&m�:�T2=�$Hb>R�>��! q��s,�ɏ�6�	��z��$'�Bh�`�}���

g�kQc�zK���r�k
��4��!�T�"c�ņ��Tf�n
���/X�-"��Rz��(
��P@�Ƶ�0��
�_��]p�Ȥ��IU%�^
}�#/�ߑ��`xur7���cEyT�� ����k��T���3:�A���_�۩��ܑN$*$���