BZh91AY&SY�C m_�Px����������`_����:��P�M4���S@P��� M10�@ �  �  ��b�LFCC �#	L�)���� � � ��b�LFCC �#	�4jl��I�i�������qtH�$� B��@�?��r0x�
�/�`@�A%���F��R�$^4(L�G{Rr �@^����4׊�7��LJ�4ˍaXV%�E�p�I�Ra�p|j6���b��"1�äMF�)�bL�y*q%8����r|[��>{��2�,h1�o ҝ�a��6Rs�C��r����A�r<�@[V�	�J��g�l\��$�fQ�,�rՌ��2���{}��4�""���F́o; �|�lN�1�歸�,�F"q�G�n��>ᥲP3��Jg
N^��h�/����Mhd2�@<��(ΎXᭋ����̋J�-��҅�OC��L$�Q`���CA
��w-	`�V����reަ��;u�MK��$T��X̂D��&�,u��q�P�\�"�Z�Y`��
)]&FbQ��@����P�c&tҌ����C�"��AE&�fei B��@KL*kzׅ�õ�4V�y�cpk����Κ>�DHBB�I$�
"!����u��$n�rɈ�O�#�#x��Q(�i��@����L�f��Q��m�!Y��s�&Q#BQ]$p�a���\�����q�= (���#�Vxx:�4���q�Te��E<���M�Fw���E5���b���|�&��E"��xG��mĈ��ͼ��Akf�c �	%�}$�ؖg���bDM ���ՠ��
a�!������oIyP�>�%�Ռ�5$2�o`I|�Pm!�̊��� �-ܒx5@�kk�cf��u߈��25*7˃UI2�����)T#�B��5"$3��\kW�����T8��#��|�;�ᴼ�TJ�O�v����@1%� ̈Y�Nh�:�m�4e�&@eT4R]�y�V���Z��ə4�����K��1%��l5/,�H�k�˹��j�bБ��^���A^���@e@��u��F�a� ��@�7=��`M	B ��ъ�	Uocc@��AA�M��F��ʓD4T>��M�M�ٽ	� ��9�0���!�������g\���qi�1:��' �$�w��C�0g?nbK`Q%3���^\v.��������Pm9�g70�bTp�4�վ8���XEo���X�BjOE���K��jZ�H� �P8P-��Ak%�RXB� ��d��\F�7�Y�I�=��hh`d��c)��$�7��|9nmx�-w�d(6уB���u?�w$S�	��10