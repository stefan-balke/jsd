BZh91AY&SY�� �߀Px���������`=���� � h��OS�=Fj h     �E  h     �eG��@  �    Jd�M"b5���@  � � �`�2��*H�hL��&�L�G�G�h ���Q���HWI�c	3�B����Wm�|-�%��O�?�U��&���L�J�*��j-d�+XҾm�ޚ��%5�O�q"�S*��\k���Eg�-��>}���f�@L�v�R$�wR��1���0�v����Nf_�7�	txC��FV2��tV����)�r(`4$�����("�D�AeN� �կf�q�&f�'���Nd�V֚�S;md�x~����� �6�8Û���l6	�|�<�0ő��̻@h���*z����A�����$��䛊�b����V( B��\�g�j�;��`�� �f"%��@�LE����Kŝ��EU�)�Y�G7U�aPk������*K�#��E����5�6�B���@B`=
���Z:��WV(,��B�0��D��� B����	�
V�U��B*��!�*�H���Qd�K��uj5�9�X�/�6k{ wk�1�
��E�HA����X����q�^h���%�u�$!-I$��D �w;h;���4� *|�9r7i�Y�"��40p�Y��-�Jjg��JC�!!!!M�	�T�e3R�i�K0��˔Z���[���3'��4#?�[�j�� �.�kaa%���2d�@��PH� \pl.x�I�lV|��ۚUV���Qi`��|�D1A�J��w�����t�_����ϥ[ԃ������^n8&�KC���O��8�O��}�O��(�؃����bb��C�~2 ��CF҃��C�e܈����e���)�����z�YƖ�W��n�1�����R%;��S_����}��e�*�{��M<d�*D�z��f��_B���6x9�3V�s$���/i�?\xp�R����:�۔wxe��]},q�*1�8חLg#�`�X;
k�uwr6���:�h4�8�,[d��5�|�,��򊍳����.h>�'�*;�{�Tq���7�f�d�%��C��J�-/Yh4���;��$,1U݆�ƈX�Q`�]�.*���T\�dB�R��'��\g(=�ؘ�ny�H�H�_����9���m�����ny�a�Q)�{��3^A]�t�(����0|w��5=o���OL�*V�S��R�T�j�u[Xl�n���˦��і����L3���%�M~�(2iu�Z��i�R���鉫MK��<�{t]�(�\�m���H��{��J���w�8�P���s[$7^,��c��eT��&9��i��hR���׎����)�5n�