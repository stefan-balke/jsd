BZh91AY&SY�� �_�Px����������`�ـ��:i@	DF��cSORi��C'���C@  ���I�dSL� �#M�L�1�2`� 4a�����44�@� �4 q�&LF& L�&@F �"Bji�S�����Sɨ� �z�@'�HQ 
������FD��4)@L&����n�1	Z4*�*� h�jR��+�}�/ݍ����v{�ۑ��ˎ8��q�q��������8�0_Ow��=�S`@���;P���]g�k=K,�kz�����$�4o��t��w����8Rb�d�(�0����r:DkJX�ޒ,� f^Ǖ�h@���e4��
�ڍx�AmӔ��W��Ɨ������1��}�å˄��V��G��\{�q(�a�=V���X��J'�T�^x�����I|B������LQ^��@�B-���rb$�p��VH��J�d"�Q#v��!jhǅ	�²�gH� �Y�讻��EUĩ���qP� ��b�.��ȓư҄�(�4QH��/�j�0@w������b�6�Vbg2FT
�����,d�F�G*ν[�Vp��"dL�uh�9U0���F+�X��4%d��.i�V�GժJ,�D쨳��э\�[�ښ��`B-��K�*t@�f��il�Pwm�ԩ�Ǵ�lcc��m�4$A\�^��!v�&9jT"�zS�)���Ȗ�@@@ �Lo�5�H�)!V��� "��fd�L)H%4�
U�ਈ�KKE�H�HC[�� c@6+���o���vby�~6�3��ߧ�ҫ��4�4��#~���DLχ��
d����L�Q�}�[�elm+b��*s���.�).f��("��aձ,�����\F	�B�y���a�.�P*����D��/A�v��¢A�	4H�<�4��f���J�L�^}<J����A"�H�y�3y�$I6�A�ބҢ�X�@�sc�PC(���bI��!�X�Y%��I}��\�p3Ϙ��[Ԑ�l ����0;�� ������F��4��/���z�`���Cc5�I�GG=���ռ�xk�,����{J-��M\L�c�ˤ.��r� �`})D
�]���[��_�ADʳR%~�H�s�`4p)�}.P�-9C)R6�A���di��,��o!$�������@�Y�DA#�E(��t��Ҋu()4T;
�"&Ȁ��y�׭	�O`$t
`3)�%H���T;���K* <)#Q�:��,��|�xе�b�{����7��Ё��2�:�#@LDϞ�iS��1 ���Ӣa��g��Z"A�1��4m��Fh5���a����ȩ<
��;����H���)���5�Y
�VԐV���%��暝PB3��0i�^�榓� ݸ���z�1�ˊ�g� �T��^F�J�Ś�"������]��B@2�`