BZh91AY&SYIX�X >_�Px���������P�]�v �]�T(4��"S)�h M  �d�50J�A�M 20	�� HHB)��h#C@4 M4�	���dɓ#	�i�F& � �$��L&&I�FSb�� #L�ͷ��-&0�<H����*���a�PЬ !
k��,p9� �C2a���:$H2�4}��nmQ�x6�ܷ5n������lWUl��%� ?������0�o1Q���u����[2�\��%U`�G+����U��x��x��e�]}���H�#)s��|�ѱ���6Mժ�f�;4�Йވ���8T���(o|���p�0cϥ���؅ĦXd$�c{�Q�����A`8G)j�W6p�F2�?�\���Z�<�L�;�e:#)�F�Ml 3	�1jƏ�jvsY�%�+Q��ݜaq��5�*gN�88V�ZA�D�j�ҧ��4����Z��Us��d�,:��6��W�0��	C�V#a]���B� Cw���S\�2GL�T��2V�R�d��h�

G�bc����-�0�0�8`�y��SJO�h�3.��%K5�� �rʐ�(I�;c��m�����7{�᤼�r�Bw��%J$���!�r(�2dm���^���ڒ61�5��tX�,�M��020���*
��%��������~��]=L�n�p��@q|Sϯ���\���qM��ơ�h�d����+��?{3r���`����+ }f=�N��������M>u �KB�9��-�r��0Q����!'���!b"i��>d��Nu�)}�8���.��KSz�ƖY�e�$�w0��g�2�s�O:��f�Z.�ͦ�5.��5'T�"�h�5�_V���Czt��~3mj��
�a����g2�+�m+��#{Ct�X�\G�9>�ٱ0b~���K������LϿ��i�*/��x�*�X�&ɡwλ��o�ξ&�s?��4j�*K-�=��*ێ8��芓T�PM��A��x��+�z*��4��݌�r�T63�Lٜ�6�ͷ6�� Z��Ab��$$#K�K����qS':׻%���$-��Wy��%pݽk�3
k|��`�|0�d}�Z�>�;]^%lzl��r�R��אɄ���Ĩ�)E<��(6�L�翞igw.�v'��2�V�S��L�/V�
ȠJ�j��VP#؃�E),�Hx9�#ԺZpR�Sr�SQ̩hqbt�gѡ��JO:�k��km��3wԍ�
��RP����7�(pL8M,dۄY˦ǳ���{\����Sk%��EDѩ�����)�J�Z�