BZh91AY&SY� ^� �߀Px���������P�q ɪhD�(P�5=������<��� h4���&L�20�&�db``$�i6��O4Ѡz�� �����&L�20�&�db``
�M#SM��2��Lihz  i��=M��/$W�BZ ��$����U��Pw�*&бf>/���w\�%�CG��:�H́���{]\yq�q��}���>��gze����;;&�Aqt鍺�n��Z��?��?�~n���o��C�v���V�[y�����5�F���W-�Ls�Ŏ1Iw�r�{��)���Uc���~<X�h`ǯG��>�1��+�ܷK1z��R�YaZ��"����y���^�a�4dr4r���_v��l����!ŝ)g�i#q�̪.;+ʪ��i�5�#wi5-���a��11�d�f�i�;bVŠ����Hl�u�a��3\�66�PͲS�7ޫ7喣́|^ۼ������������ms���������z-a�r���6�m �=>s������#�
@�=�%J$͇�`m8�Qԍ����E��(�)��Ic0D�; �ZD-�#]�~0CQ%Ҳ������ܤ����Ј<ny��>N��/ˍ���9��Hi���	�0CQ��F�O��X�Q�!�1����!:��ℸd@�*ۢ��0�m`���C�Z6n���M��%�r��v�n#�xrC6��ަ]O���Hn���\�	Lhp�eR)joS��R�;��$�5±�4�Űz4��ݼ�+".WvӓW@˜���I�`ki|EX'�;q�e>=m,�e�PU�1t�4�<���sqo6�z�f)��������e�VKB��99�]�>��nB��t1 �[C�rK�Wt���������v����՜�H�`l	��(��ή��*Re�_"�� ��h��To���=-�/�&�������h�U��l^���>Ydp\ŀ�bBB1a.�b�`��쌡���Th=MZ���kx������3�.)�՚N%�G��r=��3,<�?��<��͊�OOS����B�Fp��)G�����w�d�iu�������k1UJ���ej�yH���o�:�����"1�us��Y�%�T�ۑq��$:�n5t���k�A��qz�]
�o\ò�g�\ٸT�#7����r��n��^������ǿ�*��sLt���b��ED�&b�H�
�ՠ