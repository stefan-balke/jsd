BZh91AY&SY[�v� �߀Px����������P���8s%�&���F��&��@i�=#5� 44 ��=���  �  hh�  ��&��e35L����@ 	�9�#� �&���0F&
���S?4�	��@=C@��=F��_]K��a$4H�!^��2� �B���S^���n�a%�в̰�h�j�F�f@������>6��,���3�53�Q==?�Û煫��R��6�7Գ�N�����>���gG(�̔q��jQ�>��(E\g'zE�x۹�{��HBɢֈ�#D����K%Y�u�G
��}�,���]�m�=x}��<�=�[-�<Ե�u�J��k/S�j��2�"ѭ��}��V���j��p�Ю釡�7qE�T����(jDa5������+P�z.�k���qb�p�h@PTK1-���!@0 5�"1FNFdx�Ζ�!6"6eIzti
�m���K:��|��Sjg/}����5�󩻇�Z[�M��/��p�ɫ��s�lcc��m�4!���t/?q�P��D�D�1|Ԫ��#v�C-�EO^ <��E��8:)#�e��P5�B���5%,"� ���G�_ޖ�3�ޞ<�V���t���M��<1.g�Ϙ�k��� 5G0O PK5G���B�ALvg�Ǚ]̆9LB�*2���d�r�f=�һ��!�P ���U�=��ܘ
]=4���!~~i����$�LAI��l�oL$�8��{�ȾQ��'������=F��'��XƔk���wχ�le�t2"\�ڹ�pq.|�I2�B5�_Wa���ٝ�pg�&N^pCI9ɇV�A��^�����ZX�&	c�O��}�l�d���uळ}��y֎��ُ�g��/[<b�+_:��ń�5��i�QN_y����7�F�����\W[z��ێ8�����]�D�8wz�Q��̯��q�S��ɡn#e�U�l1���w֥�Kt�("���a�!ĝ�	�l��4�v����,`>c"	vH.�������py]	���\����=�a'A���-0���*\Y�*	M���hZ
�����=<ax���54<�CIؚ|���1UJ���Yp�|��H�� �	�/�23����F5�����-�����e�0n���7��a�*k�\:���(3������q���_B���l�Ԕ���=��C1{C9��v��wYc���U=�:pi��j��ED䔋�]��BAo��