BZh91AY&SY���o �߀Pxg����������`_y�gNJ���HP	MTzS�&�6�����h�1�44	�Q�@d     T��JzQ��      ��D�e=)��驓��=L�dd�4�dɦ�L����0Fh� I BaM4���OS&M4 &���Ȓ�䈴0��,�{=���8!� �TC�XHL����p]��B�3,"��j��%����.�������k��v\��b�r�0�ֶ6�i;�V�Gt��	���`8%d� X���Y.¿ҿ
d�c`uD��3�xDff-h1ս�\�9���Q����v�xw�6؆���ǉn;�L�э�%��%?���=l�0ѫ>I$����USCZ�⍝��ͱa�_/���z��.WX��`ǿ��u�����e�\�V��ǒ��;�����`�&�"�V�]�*5�� d+ 8����fq��d{�p��'0@����.�r��"T#Y^��me��qnb����kB՘��cY/f��A�њ��e�'�-��K��ː�M���\�f�L6(��@لOVl��I���a��Dc�%Emm(4��hwR��C-����غr��L��*�UH�e37TF�b��s*�̆NL�Y�+�&��Ϊ`b.�2]��Պ6\��J�|͊D5��kA�-u$;3
]���e%�UW1t���x'.���!�1YXRi�����S�/V3�k�"��ՠ��Qm�*�t�]��)�Q<F�g�1�RȳF;&��T3�����K\���:F�61���CI
�����#�
;��%J$��!MƔMFF�EV{�R���$FGMP�k�82�!��D�	MT�_V�5��-�

��g���&a bT��z_����DF[{�>pd�*}��q�F��qn��s5B�nS�y`�Xђ*$Jj�+��pI�<*{�&�s�䙎_b'�q�IN�K�<�G)"z�׃��<���oY���RD��BƳ��C�ݧj`p)hX��̅����M-�d�H��=)�)����Jp��Q�{s0�"������R�;�<i'��Xƚ�0��M�ANG���Ѩ�KE�����w*��LNT9J�)wyk/��>�xq���L��_Q��ʢ�RIV����dc�WC�6Ӣ󝙲^�0]�}�w���K�;���E��]����|��/
���b�M���^-�,'I�_=+�e4|uo9��[~g>��L�R*�vO��\��e����I�k��G�����G[�j��������CK�5!}�1�p��R��PX��l:$#H?"]"�V0C�����\Tу��Ik�Epؓ��J۝�Б;]I0��HйiK���f=ۦ����s�㉭Ǻ�v�U�̻��#2�"u�C`TS�4�(��t�N��/|:&�Nׁ�l.{����i�@Ξ��1�v9�DX|�5�۩���ujLm�:�$����K�/�V}�$LZ.Ye����s*Y.���19dgљq�2�����z�e
9����˼5#gƸlo�(�:�=��z��.d�41��.�8���檘����l�4�ش6���ڙ��w$S�	�:��