BZh91AY&SY��W3 �_�Px����������P�kݜ���M�%)�T��LH4�=F�&�  ��MI� 4      ��d�4�����T���4��2 <�0`��`ѐ��&��D�!'�*��4�L��&S�'�H�CMf���'�HPI@�����to��ڀ���S^���$p<,����fA4w5TH�F$Ϸ�ǳ�Ex�~�����K�M&��S(�?�A˔�����G��	,�~�pJ+�цw�99�}V*�`��;m5Ԇ��n���p/jؗ���ks��BT��I
�Y��#�P2Ã�J:
,$&����NvKPAQAE���hs(]W���數׉wb��-R�^��y��"�i�U{�`�E�������!3d�dhBE�FE5�'Հe�X5����#��ROK8�I.�73:�8�B4UJ�� ����Zg����*��zY��q�V1[�߃!�%��U�b��,�3ȵ��(���J*&�r*D��ՑfTM���z��F�a�6Z���
%b�G���61���m���y�t��U���T(C�y�(��HdSoơvK���FfA��ے��h��DS��d�+2ʠn�B�Ҡ�a�՞�������람��g�|b�Aߓ�қ�p�$��&��٫��E���r����7�n�H��(��|ļb�G���؉�L%�;�3? �������zõ"�B?���1�Ȇ~9]�S��AB�?���"yt��̴IMLGz�Ѱ4aԠ��L+J�s��,B�!�J���A�,�$�UJYmt����5L�DΫj���2`������r��&W�����W���0l�w�'\���X�@��r%�
B��Wa����,B8q��I}�H�]4�x�H�gD4]T��~|�[��%�H�j������Fr�֚t�Q��/���Z���P�7!��*h�xu�p:	�Ψ�L��4cY ��JFHnW��(h�(��As"�|d:$#H���D�Д������Bb���ȭ$D��F�؋z��	�L��'H`^��<�P;�ͫ�v"@t� ���˺����2���u�
bPh`�gn�F1>�+Jϴ�,ax�ea�XV6��3��eC��1��0A������W�W���㠸qF\,���k�]���g��6�PU��.���:�-w�Pg��v�:�aR�V����W�4���7�ZL��Q�BAkA���̖��Ԉ4���isk�nT��}��h24-Z�?�w$S�	
��s0