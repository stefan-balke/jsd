BZh91AY&SY;�� �߀Px���������P~p��;q��0�&i��ѐ f�d� PS�LMF !��F  ��$�I����&�z��� ��& �4d40	�10T� �4�&4���j4��2'��Ʃ���]$%�aĖB��䫶��ʢ]A��O���UU���U� q
�Ħ�\�`���Ύ֍kf�z����W�Q#���V5�]��
��J�D�rY��ԼR�%o��2��A���}��!R�c��=&Rr��R��%����(�Z�4h�0�����2ݢֶ۳��l:�,��*QJ����{���3Bu��yǷ��e*�|w�L��G��H�����qc� �Q
���%�/V��Q�(�t��94���LE��I�ʈŰq`�29��)�9\h��鋍<`��O#%�'i��R�$׺����G��{���
�����U,C������luX�J"���`��ќ*�HBY�I%�3w!��<ʹj��$���Z��Щ*f��XB�GM-Z1��-�$�11��r�DPCA�bL$��@�q�G!(�t�җ�(�J/)�#� �NA�2�D+L��uVf����r��n �Fy��$��̏�گΊ���;�g��I���u��!�9����O�}-�;ѣ�H~šcq�竽n�}I��)hm���0���L�$�^�2jX�NO�&)Nt9O�sDh�*M�c:�DB�P�Z��E�+�O���gigZ1_�U�T��:Rx�HQ����[8�|��l�&#�iy�0GuBUUUJ�V����fe�W�n+��G���X�~���ߞ;��)�+�:�۔y��{{,��8��bq�W�3��0}��5xm�u�>m�mqCN�ƑbŵϯR��]���d�RI՗4=���*<l��z*�8��S~�k�C%�6�]���Xo������a&��d�gA���Y�M�E�;hV2a���L����8I�zD�]_G$=��z��f��R</�4�{�������6��W�ਔǹ�x�א� �
��y}]ho.���Y��KA�O6&�T�P�oj�R���׌mh���)˟M���-F�Rmt����"���Wk2j�֪��M�a�R����F���y��o�B�/�K��F�
置��r�/s���(]�����vt��鮪|��T�R�"�e�
�F&�e�.�p� v	�v