BZh91AY&SY6E �߀py���������`?y�[vq�  e� � J24S��@ h    �&RJ=@  �   ��4�	��0#F�` A&�Dҙ0F�h Ѡ  @2d�L&F@��M#4i���$ƅ<&S ��jx�`����L�$�}�dB]):���Z�A�q���vO�f2K��L,CB}��5��TMHT�d�e�J3 �`�u�B�
�k{=]���z����iJ.%):N���n����|9�ɍ�޺��]:~��aY\s���:b�Vs[���m��X�7�����f{ʙ�T�PjJ�SS5Q��Ä�a�tA-�4�ph��,A$�R��f[j�pI�s{x���3M[Md��hcf�o�Vgrno;Nw�$�V�ע��c�#�'*�UUTTD�Q�k.��s+|f�!|!	�Vc�uǹ0\ ������@���P�u�Y^@���;�{�W�����.ԡ�K7�5�,�C�����`l�
X,�� �0#��$ %�7!4PA���=�?7�A�^�*���Q�0�%�+L��ڪ�Q��vu��g-ñ/��X���M%�	q��8�w4���<Qp�����k���@��X[l!y h-E�$Ag4�#LY��Ȓy���� >��=�bES�X(���rhl��S��j&Y��*�ڙ��r4=
��!�M
S�)W$VP�v�|�[�oIps6�\D`�Q]㨹~\,�6I��A�ܻ��sԡ�@�y\�n�4�t A<��B�	�m6��Lv�a�Ļ�Z2vEN��X9���x��� D��\���\��yīE�1=��]a��a�������x����~�]r�uQ�����US��U�4S��ʙ+�(��g��<�QE�Ub���8{'l�E�i�(h�,�r+�ʺ,��U25R.FbƩe1`�cuƖ1r�SE:��Y�P�U*8�B��(`�QL1bŀu�`�t�@�Yp�B���&��!���*�Zg�O��o�"�����Lq���R���	�v^N|OHUr�2���$�:�/���k�TG9�z�Ņ��(�㣴zd�d79���#"��؝;9;��>}��$h��KH�����[�ok�/=)KC;��u�H��ĩ�\�j�TeJ��I�@�F�p?�S����_*E�	�稜{�;Ь�.��6�*Eh���.�T�����`��ҳ��)���I�R
vH����s�.�oZ�,u�VS��d�u=ZJ��$U�X<;̌|��֊������7��{%��?���������q�q�&�c��b���{�C��s�BTeu�NJ���a:ͥ�K݅M?�yF��h�7�9�$X�ms��ԭر���9IRg6T�oǭ�;�2*<L^e=F���6�e.��2X�X'���E0��4Z�뭹|Df�,]87���C�u���(d������3A/§B�}�+�ʌL��Z�Zŵsn���I+�;�B�S7ќ�r��ے},�-ibx�K9qS���r���I)�k�s2] W�Fq��JN��(K�/z�ΦG��4'l4x�Mf
�W§N��*#
�\��iD��g3%7��62]k9�Hf�̗�/�V�] b��ׁK���=���K�l�bӭ��&���FY)#���U��L7ݜ���f�񮽭�%"{e�����h�R.d�ic$n]%��X��j�=γ�~Tک�T��Msѣ�]��B@8�`