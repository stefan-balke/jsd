BZh91AY&SY�ط� �߀Px����������`~y�6�Ml<�pX��2OS�6��   4  �4!�I� h @  � �&L��L �0L�0�BEO��MF@yO(��@ � �Jz���ChI�A�mG�� ����	Ђ6�УaO)��d�  Ѧ�Ҡ�� E���B~�Y��(��4;�D��,��m��d$dhXI�a4vڪ�)$���ս�c�ٲ�:��4�2e�0�ݶ�BՈ`�s<���4�mB#�!�Ikq�P]��[m\K�x9��Ӥ?��eFX��s��A�jqF[ILKI�+?��'�4��ƔHK�K)1����D�5�I��Ȗr�v]f�Hd��`ņ�,80Q!� �r�Q�&�Y�[���{ٜT�"�9P����&,YdN���tT3����!@)�;t(b����4z�C$�'����;̲��v�J�&DM-'!V�X{�<0�ĂY�/X�5Db�)Ţ���R�(�a�ivfg�`k(h�mWp��&C$� ͔Y4dpV����iZ� �FrU��_M�/E�S54���E4)٘�J)ub��b�	&�R'ZQ*�jԝ�RRY�O����!Ȍ�̑z��vyc�-��h`!�c��J���T(I�q�*Q%���	/J�/��X KX�S!�$nH�hX�A�j�-T���5j��-�J���kwR�li$�E���m�s��&#��� �~6�V=%ьH%��A�2lh$B���aD8���%}W.��hl��*Ͳ���ֽ��.,w��$2 @q���>��N�ԯc�E_�Q
�i�Ό��#h`����Z�~]�ŭ�Ǭ�j�1�ьE�*�J�-�N��{F+"B���WB�!��}C��� �L3I=�Pk���������Ph�DP��\���(%�1�"	u`�1JR�6u�$8��,jW�� �aD����_�������j��%�z���i�{TI.��1��v��8#��o�4�H��iT4g:!h�4�QpJk�L�c�j�{�s�ٙ̒\q�s���}K߸3U�u��K\ ��#�zIz��:Jz���@���#���m%9�Xnz��$$�R� $j�PE�;�âB4���H�d+q��R����6��.�"l��~E�jΌ�av�]'lmE
M����|�p�Ҁr衘о!��k��w�����cY� �ŉ�!xՂ��Qj�+�;N� �cK��|£i�::HcH��m&��S���ƴ-�c�Q�p�U�W刲9ZE��&��ID����A�ff@���R]��	c���1.��,Q�unB�R��Z�_�ay�, �(g�7��X�bU%�H�����M���ka�3���I�B�Y��.�p�!ͱo�