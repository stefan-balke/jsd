BZh91AY&SYh��v �_�Px���������P�v�H�� p�4��OJ<D��i� �FF�`LM&L�LM2100	L�MFC@Ğ���4`�F���a2dɑ��4�# C � �A4�S�z�� 6��ShO�BH(�V$ /��9��*Ф1$��]�m��pЬc�Тdm X�^Y�y�j��\��]������w����&�Ǥmb�"ĳ�[�wr�'Ju��L�̰e�������39dj4�\�]��ݢ3Z�O��o�H�>+�~� eʜ{奥��1ݟ�!���l�Z��%{)5��I|tP����z3�tr�V��b�GO�An�~(T�;��a�M�Wo�D5DZ���BV&Ƞ�QpP�����@RIEY�XIZ]R�l��BU����R�ल��&I�c�����I$�
�Ѻb��ro9d«ߑˑ�ʰ���%"JҖ	�m!jjEQt1겗���@ڿ�s41�a{>Q�����k�[fw�k<�BeD5Fܚ�h����b�"���z�-
q��@��S~�1�:�Gy����
fb�����;%���C����-�`|@fkH����)��+ >+���}F`w�pIxv�d0���l�}�9/��SD3q@�y�2�ēʁ*��i�����Q�cPmd"����3TL�ޘ��&P�U�)T�o1��P�d�K�݄!�48С�y�->��0{���)��I�8óʸp�\�$l�Lg&vA��s�-���ڡ����۷yE�2S=��`e�9m>Ś�f&�-�ka�`^=+Z��܆�FKF�k�x{8�z���m�^y2�pED���3PV�s���(�/ d��B�nPR64d�B��Sg �9�&�h�P�"&��F�'�V�:�y�@���	G����ߙ��?�ǣ������XЙ_!�s��>�3M�tv�@��ᢸ��:�C�^Z��ӽ9yFHcUy�"cX�[�A�7p�U�V��~g$XN�5'u�� �|�3i��0�^5�T8T����t���Q��NƑ��ߙ����p�6��"�j��g$��������T�����j!уB�#��3rE8P�h��v