BZh91AY&SY1�� �߀Py���������P�q��!�-�L�	$HȦi��?Tz��� h4Pj12��L41i��M0&!�0�ȅ=S��di�z�    2dɈ��	�����$�&�I�Oҙ�zjzL�4 �6�'�ּJ�D�����.B��ߢ�lC�hcQ.���K.��?�*���J�#(;j&A����WW������%�wn���x���:�ĢG����8��ek�EkE)BJks]���Ջ�~�9߄�x�7tޓ0R^45�<�2b�%��X�l<�,Rj��&����Bbb����Ҫ��s�̾Tuѿ�2��L�0�Ɇ�7�`o�r)UR,���#�m�P������}�THZ�N?h���h�r�zV�"T\D��r ���hM�eڬ&SVŶ��
Uq�"����mM���j�l����&%(���Y���/�&8Bla�dQ���#':�"��1����A��Q��Q ecF|�IS"
���0�{W3��:')�$!!	m��J1�����ܘ�^1�,��gڑˑ����%�Cw%���.���CIM\Cj�#b(E�2�̄���Ds�ə!���`���ۨ��Q=�tf2�ά���X�GU�i�L���%u�օwr��(�؎*��ۓaS.s_9փ3%�>P���U��zϔh�u-!����3[��,�r�����.��k�o�{��|��>謕A��x�%9�"�Y��<��%�jm`}��Ygz~��[|�ODIP�g<5^4�`Ñ91�=��E�7a���pP(���&�8n�e<:Y8��ز)%[���F>u}c`li�W�_�"xLC#pv}c}遒g��m->E����c�4m޽nlb��l"m��,4��r����������.���UV�X-�x�5+�q��䊓�l�sc�C��w
�+�vU��N=��oLT6/8�_F��J�r��@0Iî�V�����=C�A`�MѼ"L�r�j1=,b-}-bڞN3Ѻ%sa�!�����m�q~�Å%�%���_�惼m.�r�Y]f�D�>WS���3[�l���R�qy�Hda%���3hu�N�����0UJ���\�Q�K]��v�5�Js��1�c����̗�_,��s�c!�;�Yk9�R��=ui�{#�Y��q�B��`��OO��$�	�2E�[E�,� �8��3�M�\ɶ�f�q�n�c�~���n�e����A�`d*l<�G�.�p� b=_