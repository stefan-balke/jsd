BZh91AY&SY�5�� �߀Px����������P��-n�p�2ha$��2m#z�ji��F�(4�A�A�2b��@�  @  &����z��   9�#� �&���0F&
�A&��P�S�S��<��z� �4�M+�J�$KAD��,�{}ߢ�j�~��Aa!��֛�9,4J,Hdmd�f<�����T�k��ܭ��W���U�|X�_p%�Q>���8rZ<�[u�*���Us[g/u���~����7���z��`̴j���gMA����]H��Vq
�Qi�u}�fѧ>	3��2ΙdΥk��Nq����:wIs��n;=n��
3�Y�a_\t��Q��UK�J)�v��3���Q�
�/F�����&��V�V��d`��C��1�`j����A���i��x`�'elHdԩx�J��qd)�77������tH0�QV����P���DALw��ޢ�X�CHQdJ!�uP��C�L�+�
s()��gz�Dˈt�
�%Mq6)����՗5*^�E�ʱ����t��61����CI�r��X6и��*��;�J�Ie��dJ�GR��d,A�"6I�k�*��c�1����eF]-�((F�͏�0M�6�_$�M�}N�8��+��l��1������8���r�Hv�1&~�`g�,�NC��T؅��6�ӽA�x����'Z������\�e$}��F����y��;���#�Z6]���q��L�Z����{���wH�
�y$y��R�O~&2|�Y�C)����Z�>�o�,���ڒm�3ͥE�17$`xk/$���@ƺ��;�2�ѵ4���!�Z��d2yYÖ�83��fr���m6��9�\���fo�]�a\�:��v��X�wk�������$t��ʔ�v.�|������ܹgԴj�!,[f�"
!ER������Y�J���	�i`Np7*�^�tcu`�uk���FI\��Q��Z�*�X��e�d`��K�TK�p�ڪ��֥�7����|XtHF�K�\4
ɔtQU��X%��,�Z�Q\�0��\[}	Mм~K65��#����z�2��ß�̚\����mTL�;�]���"��QM%�t;rH�_"��l���y�ݍJzq4g0UJ�
oޥ�S���֋ձ'�n`�\���6�s��Cc~k���_.��9�$bТCx�7`�5�.r3�04��p}���E7(md�w6��L��e�^�	$`�"%�uHy����/�ġ)O�ƃ�hd��i�����"�(H~��E�