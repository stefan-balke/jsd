BZh91AY&SY�C�� �߀Px����������P��v�T��viF��#����!�&�4ɦM�@�
��� 4  ����I�=&�)�!�=M @m&�� �`�2��H��#LL�OST��S�~����z�@24�LJ$��H!T�	@��n��L��Af� �( d��~hہtP �hU*ah��0�*���p��⮎��܎q_�]��Y$~����e��E�*፷����� �ۇ�Y�f�9��ˉ3�N�V��[B�y��Ae��A�`�r�W�h�!PZ�7�:{8��T���g���;����\b6�Y{c�6���f�m��0c���Z�[�i�&W�����\�1n2B��j�uc��bVb�iP��s��q���M,\	����1|�|���4�rRh���+{R֌^�a��z�E�Q!���ښ�KFM���<PMT-�W�@D�'�����Y�k���P�a�\�~�33�v�m��A⡧�5H���M�@���%��~&1$n4�ܥ��\�E-U�G#*5Y��Q.�! �׋;	�Fݑ�����m�k�?:�� 0
#L�.�v.��$1U�<U [�k���{�d���<*m� ��i����Om1H<�C�b���=��EyA� ��5�o�}�[���!�^��K/R�˙%�H>��3#�0�Ĺ��*A!���by�=̂�_jI�0��k��I��v4�X��5L�DΝth��2b4L�
	�!�XEm
l���-���.3����m��М^Mp�*
{���!`V^�(	�!.G�=�8K �71�]e�R8�����M���-��a�I}�� �^�2�V��1sYjň�p�y�ǃ)�Sv{�ű]8I-��<>��������aa�
��Jca ����nWI�P�0P��(!B[�9"b=�AT�m�qn3L����	�C���gz;�Bx�h���$6�fPBG���`y^f�D���xv�4^i�1���ʺ�X\J@��F ��G�H�@Q��6QY�ub��HYhR6��3M
#���!���1�g��S���R.4����
)wᨨ��ۂ���1�K\!HsԬ�Y@WX�qnaz/��	�0�c(�iz=���G��M�cA�

�֢�P�4��f��_z�����^bB0d(���]��BC��