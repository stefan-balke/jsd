BZh91AY&SY��y) -_�py���������`��#l`9�� QMOT���)���$��A��FCC���S���F�     2i�# `F&��4� �S$�2mD�i��dфmC&CMCdɦ�L����0Fh� �L�ji��'�~��"<�T�  ��OMOI���o�p�TPA0�����̕7��J!x�D��"��~e(x(�dG�0(�OlkQ�Q@�;��G��OwO�ù7�'�3rm��I5v�o!p��u�f�2��bM���,lR'�{��p�՞T\DQ	)ǋ��%�2q�+�n�Qc��Ke>������NYi��.fjL7�n���Ү��Z��w^_p�]�d�r۳KX@1#5`�J3-�X.���)JI�V�o����q��,�`Bl�����D��]v]��>Dk���s�5զCC�E�]�[�7q�5���/�t�Ե��]�H�m��\�N�³꘨cesr��8j��.�����T���nN;��8�ҨC�>0*���2��I�EhG"[-�%����MḚ�u����lx˺{�U)&j������NI�H�ۃj޵��Fڒ�-��ZPN..Hv�q9�����|��⫌P̂a�U�ґO����HT((�@H��4J�@W���KK�U{�Ӽ񝅄w���ae1l؉U�W����.�U���Ue��QdE�q�R��
��"9M� �Z#)!�](Ct��y�j��fooZ�� �ED2�������L6�i�l�`�-D	�"���"�WK1�R��_J��7���:�B�2I$�EUS����Uts�82B�߃���E�-��D��H�B��T�T�%IRG��*J�����Ё�1P�l�I!l��"��UGmE���{J @@�v���(�!"�U��C$_�T�zK[�`�+�2y�ڧ��0��܌C����C�Dx�϶g��*���=�~�N�$����R��^�^��g٩��&.�*_ ����>���� ��e�_�B@�<��H�"V49AF A�gM3���C�~����+c�É��\a� ��lG,)����
<̼U�
��g�]�� C()��Ӱ�ѡ�
%���N��R5�̀�� ������O�=ؒ�>}�&�?[D��H))���ds�>$����M�Pjfj�h+�=����unP(��`J�S�ӿ��2��`Q8]"Z� ���zK��["�*,@����!7���@�^znz���M�ר6[��=�is�B�E;Q_��%���@�`���k���恑 ԰o��`p�L:p�6��C�a��D�N��ƪ�􏼺�aȆD��	H����L!J6��W����_Q�W !���(Ԃ~u���噸�m
����`q;�X:��OPp"0���9%E]y^�5D�=!@����"��ŏ�K���z�f���V�ch\��B�HT���`Jh!��������oD���EzX����Y���"�4�	BP�mv��4C��v�2�"��$�-]�еkt(���_�)��ξ��X�==� ��)S�h]S}R�gm�v�#�v6�/��C�#��ם����)����H