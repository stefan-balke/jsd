BZh91AY&SY(5� �_�Py���������`}�@yy� 9� ԓmSOH�yM �� �  �O�FD��Ɉ���`LC F�dɦ�L����0Fh� 	L�
�z�G��S 4z�@d "�!��##�4� 4 @E�i�)�2l��Mj4����$��e@���B1|v�3%�����@��j""A��R�hUV;��H2B
�k��;��W��;�}h�ޗ������k���*�Y|Yyv�l�K�tW;�KK9Dc�he
��Q�#)�E���'7���?�_~ȔR�1�������|r$c��1����x;d��,����yj�D�1�cn��Δ�)"RnR�(Z_��K?q0� Lm�<s�����pn9��U���}�8�M�ܧ)��Nʊ��*R��C���T�c��M��cʨx�؀�����TQlD�ج�ۆ!��F0�Ѿ,@w��,L������+�#�`��i:�dZNB^�j��x{��aS%mN�f���B����Elrb�Wrb�F�p�m�����#BTY�NL�re�2�n3�fu�ad��XU�hY�(cy�UMK%Yˊ,��Ä�ppUI�Tr�ҺH��S(�t'�NQ���;s����VB�hr6;���h�*�br9�5%b���6� �D熠�9��_ �aC�D����~lQ0��!� ��x&thc���&��s��d�g.���os3&�ż����=�!	K�$�P(�{�_����r��~G.F�݊2()D���!:�Si��HB��!!!! JD'�`���BBB�pG�CA�"V$��0�^e~���6�＄_��U����m��o�p!ɿ�j6 \)#�U-� {��@�<2��N��#0�'���ԅ���`b"#�QD��s�D^/�a@b�����p�J�@~Km��e� �	! �,��[�l{���M
f��h2��Ac9_���C� ���5>	������`�3Ba����W�$�J��x�`�csy��Z�� ���]LɈ�Mg@�Ws�`�R�t�bx����{Q!�9����^��@b}چt�Jb�P�i���<�L�m"�ȣ��ʞ��n�D(���HZ>�5&��F�e�9���3�� �شhז�p�)ٻT4lX4$���w�0<��[&�,J����Đ`�)H�)唣I$��$�zp�$(b�xI�X��}�f"�u���P`4`��H���B�/#?w R�J�AI�J,���Ǿ����l�適��7%����A�2��9�"�W�G c;7 *��R<�V�<��X��a�$4ӹ8�"@��B(��r~�p(3Mx`*A�8\$bH�Y'P����$�b�@fF��l��+m�B���rF*%0���G�G��c�{�5i1��˨�-`mr$Xj�*�g@���㱵�pS���f4F
݇e���ܑN$
A% 