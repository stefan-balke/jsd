BZh91AY&SY軂� 2_�Px����������P�]��Bp�ѐ+	DM��'�yF� Ph�2 5=b�C4ɦ ��Ѡ���S)�@�����4�'��z�db4��1�& �4d40	�10T�&LL�e2�I�Ѝ0�  �m'"��p���&D�DY
�{�5\�tA��I�� E
k�{�ۂ��\I�%�
GST�H�i j�9�&�>^n7>����4��6�E����hT)
���|m����P-��t��X��t�֭�H�=qH;��و�RX��1I���4�L������1��3]h�/�fӚ��&'|l���(����;m��:��H ��c۷�!����b�i����Y���Ym%TzVҽ�%QS�~�c�u�V���� ԝ�K��u��^鴂�P�!�Me�a��L�c4f�"M�!�������.�)��a�K��(�ki��Z'��^г�&+���>R�=AĚ@�|Q���i��@�҅Ȇ։q�x61�U8z�|;�2�X$��BQY�(\�L&�R,E-=�CQ���|��x�T��^CFE�a��3f�3c{jT!���g6��YV�Ga�61���m�� �<�<=A�л:��B�w�z%J$��F+���Չ \�E�������2�oG(��`�vPժ��[PP0�r������&�0ƯK/||��]�#z��3N̾>�����	rE]�a~�Ǚ�q ����:���h�\�8�]�R�Z�u�>�K�F?e�cl�����;}���Ӻ��,r��y�v�<Ɂ�Rа�gϐ_��|T��$���|�U9�$��g��JZ�]����Yg���$�\cׯly`q�<\cѨw�.y8����ˡ"b9�+�C���`�����8�í�T��ʩUT�UTJ��1��j�C��|��c3��\b������c������J�r�O����x�7�.Y���B9�w�rZ$Iy���{o�J��X3��b�[U߸ҭ�e��x�	rk�2�H݀=^G�Tu0�+�WX݁��Y���^��y��}�6����ҺI
9��"�%�3q�!̗H�`+�A�Y[�M�A,�l��O7<J��h<N1x����T������jn�ƨ�x~�7��;x+�ڨ���y�S%�+�r��(�K��f�~��������I��#F�T�!N<,P�նZ�z�1k����N~�ړF::#��+�/ľ]Y�o`Z.R�S{KIȩd��Cc�F�Y(3�����v�X@Â��5>�o��p���m�%#ֳ��s��P�/d�41�-�eհ2�2�g-GI#�<E@�PT��.�p�!�wP