BZh91AY&SYZY� �߀Px���������`?���A�   %Ti����@  �   ��%��@     sbh0�2d��`�i���!�JzP�        ���&L�20�&�db``$#@��=G�e0L�h�bLBO���B(	�����#2H>���
C@��&I���m��@�
�,��Ƥ�I+D�#�N\W����z|G0�����9��;ٶve�vM��vL]�0N�ɒ#��@�}W�\ xf�褆ّ)2Á���2��,�h����Az��M_!���s�2�,P�9�0���X�2y�H2�H�NR��\]>�֗��4�H��Ә�U$�!��J�,��"4�I�h��]�����t�	�y��zC���h4f�[iN��8̍s$�8k�E�AI��Z>	Pb-j�Aȉ5�����\qR�6�dȁ")ݭhDZSa�j�2���ԇ1�^���g��e�	�:D�A@����f�32���tp�$V�RC:���J6�8F����	q�6ܔXM�k/��ͥV��c\]�H��B��+]omM�J�՘+L���W$DM�����WW��Z!��Jڭ�2�5�Jh�H^����Ď.�(��;��f��b�!4�h�GBLS���M�4);2H*�SW�1Vd(-E�ў�S@�
ӂ�r�,Lɹ{vD�Q�@�\8A��\�`-Y�h�C-i��n��H7P|�R+��UZ��^R���&]7M��'��l�gY��;�4QE�*�BUvz�?��Uw�DbB���X��$ů�\������Zd��t����-]#"�F
"��,��DB

-*�iEuR�D6��D�@��b��4!6�k�ɿdz.Lu�f���@�h�2C�C6��

��ܛ%���ѓ�.�M�;B�E�>ś���UX|)I�-�E�r�BkKP����2��}ݫ���{�ʐ]�4!{�@d�o�Վ�L;���<��_lD�W�g���K��d�zP��,�}h7�6������f��>%��O=U���
�6����N#�(5�B\��-P@�!D�&s��5�R��R�^�tZhp3�ȱ�_��6�	8�P��
���@�_�4��UE0�.����M:S�/$�a%�IU�+�l�L�]P�IM[�׸���΃�P�c�˛pg��lՑ�W�[A�����W���8oCFu���B�����W�[a����,hȸ��D�;H9�B��4NQ�0@b@9�� ��bdACH?r(�@�%Voa�eI�*�RB���ݠ�ބ��Ԅ.��`39�Β$1iz����0@N�6�(������4&W��q�$�C\��{P��& ��^X�u8�h�ci���x���*8D�0��#6��\3f�fa�8`��i'P���%�S	��̳#P�q@�B��$��%%�2�T$#ԩ�4���vF֓=D&����A"�ŁT�B� ��D�����ީu��r4��`��a�뾟���)��"�