BZh91AY&SY�H(A �߀Px���������P��ګ�g�S-@�E0��mS�����4��H h@�J4��H��@    	�5OSmH�=A�@   �F�UM  �� �@�$�	��I�<���=OP=@ h4���Q$(@"�H� �ۻ�9��[���P��k���m��X2��Gf��W���;���O��gAy�D>�T�V�@����C��Y���1Cs�,m�q��������=��q6�z(��b:�ZArx���љJ�6�.��е<�IhƂ�$+��9�H�%�L.���&�?$紘t`�v^���j��m����e�TRq�Sm�!ZTE2 �����&TAeo1����@��V�c����l�U/�E���\"]5�O�m[E*Q���,e�4Y�(k��	ȑg5h-�\*��R/,�s��%��l�:y�Ҷ�ё$���b-�Ӷ,�9x)�$S�� R�j���Z�eF�jʹ�B���NV����lcc���hi">�P�^|�w&�����5X�.�ØՉӠmL�*�扵�IÂH��L�4��(e��bI	�gK60Li
�}M��_�]<���j�7%������M|���]��3wĜ�>�}aDƼ�ǌ�:�V�r��U�T6��1z�I�E��H�B�6�]~��c�;��ć�P^x�#]��P3� `��C��%��5Oi�@b)#�f�f��͌k�I�d3�X=>A���I�J���EDݍ#i�߬���622\�榐ɤZ��4��DT]�)P�Fr��p3��VhV��M6�li'I�2	�^qH-���T8�H#Q��P��$ ���A���$�4G:y�o* ʈh��BT�*�"D����(�/���g���=60P���Ǫ��m١�BŤT�$|�τ�E;��l2�\s8���AA��Pp0UG^��cQHA�� $��!D׊"�/�H�dvl��)�@�� ��D^g�/�r�zďzU ��^ �D4��3Ȕ ŵ��%�ĉ�\���������pXI$p!��CG cq��$j	�2�ߩZVt<
��+��ס@�Hc&��$T8�F�yA�3�x������YVea5S��Ċ�@���sM����C�C�b��2:Gy9c9�a��դh��z�&��s�kX!H�ʦ\P�"�@{�X��L���f���`Э��d��w$S�		$��