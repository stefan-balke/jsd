BZh91AY&SYe�� �߀Py���������P���0ڠM�	H�MOi=ڇ�=M��4b 8ɓ&# &L �# C ��U?I2h �L���  b �&L��L �0L�0�Eb�BmM�MM�4�OP ��)�9���]"H.�YH ���{�Fȿq&�`Mr��g	8�$h4,�e�h�j����G����ڛZ���n�!~gN���h�tV�`GX�|�1��H�L��?���ͦp&2����}�K�Ć��M�d9{Db�=nRI���9�*�Qh;Z~.��O�[�a�6�������"�`�C�n�REǴ��"�~VY��1Qlvs��.&;��{�lck	f���֗�R嘲f ��a�PL�����M]Y$�]L�e��b4�4t8j�g6�vYZj��u�cux��lcc�m���B=��ऻ|r�@�8h�(���2�936��T�˓%�yM�H�dUJ������k{a�E )BK�U��~�]͋�ln�d�WD���vHS�����\4��z
�Rg&R_���bF����1Q|��r�<P�@�4ؖe��$8�4��	L-h�^$F� ��6 <��ϊ��,�����j����LL�:��)�gH�y�YxL�$��±��3c�^E�Z�� ���t4j`ɋjf�
�X�/���f�6����ei�@��4�}c���[��9�L�� ���˾yd�08�m$�DQ�T|�T���$@Έh�d����q5�5�G@2�My��Ey�f�`[�lh�@!Ҽ�Ǖ)M7�CG1�ɡ+�ޣ�G����g0��:��"�05�M���
Ź�+�Gi"D �F��d�\��6��QT]"�Z��3�K�.��s!� �fHJ����*�<�	[ P�� ,�X��2�4:�07�" t{�m7��N��f4*�+�u���PP�0���8�n� �犴���,�^[¡t��i�8p"@(𴄑1���o��3��R�����RT	(�nИ:���5�a�j�k�@҅��D+Q�"q�
hew(�4�=>�qNF����"T�\QE9�@;��mx��b���Ă��v��l��w$S�	 �[ް