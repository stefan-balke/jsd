BZh91AY&SY�x�� �߀Px����������`���u@�
 $����jy���d�4�4� M�
J  �  �  s F	�0M`�L%OҒi        �& �4d40	�10��h�zM4L��6� h�4���N���@A �,$�����G&�#�,Ф"� d�����<h�,���4w52� B� 0}��]:Jq���S�w���qJ�.a��8s��������ttE�/�������{"�J�eM�]._X�(ʪ�P?����"sz`~��a!����e��$��u�6�b�Rԝ�E�(��l\O'��
�	��� �?�+�����.��E7��5��&B�}��cQ"�,���6ҬV�����+�nD������wS�F��	���+Z�:�c}u��G����4��A��e��w4�+	�����CI��j��L�%�E��(��m5�C��2aB>ChP�ҔB,��X(�c2
��1:�ٍU%WRd�P5K:��e�G"��}S�pMX�ԥ�!�ռ�!�ƣh)��H���֫�U�aL BM�dfuY�kBP0�E[�Ѡ0t�R����D���1���)UN1�>�{��	�r��]�n5��sa���l��)	(Ø�� �^���Ep�U��Bٰ��ʔ��#+
УrmT��$��mm�+%Q��iF"�$d_z��$D��.�AT��Z\�d�T�J���(R�!����4!�c��K~_t{���Lt����9�����.a�I-�M�N{�/���Xl�enc��Us+�?�{nm��ĶȖ�4}��Z:B�
�,Y��Ik@d�H�A�A�dy�#��-@�BH+�wJ���K˹��RH8#6n>U
�����≤2�P�w2<K��O]Bmk��Y�hw�.#����4d"*uc<�*���s&!2y�0jf��6���ڐ�gǨ�ְ��CBq��`��40���@x2�/�ӄЁ�fP��P�I=W��sY{����(@idT�9���MDJ��9X8�$�6�]#�b�H.J�`�j^Z#΅����ђ�����A��;�h�-�?3�*�ΐۙ�M,06lJ�6���gLJN��B�@s�P"B���AK�"J�T0
Q��H/VZ����c�4W"�ZA�oPDpF8h�N���Y0@�8��dz8�6�	��������M �v�0�,��a�/�I�P�*6�(��2F4��D�1�|p,3N>
Ћb1A��t��QK�R� ���@hd�CP�y��p�_��������%�0��m�G�FW��g�{s8�M%� ��74).8�%��J ��ᦦ׉ȫu��fhB0hXdv�_�]��BB���