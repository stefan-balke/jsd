BZh91AY&SY��*) ߀px����������Ps�e����$PS�4��ji�䞘���j`&�0���FD�P  �  @!"j��S��jhmF@��  �L�1�2`� 4a�)�4�3Q�?SS��4��ɐ��D�сD���B*�-B @����b/� �@�!���?ɶ�;��hV���&��U1$Ϸ�ov������,�|�9�e��p�k�,>�E�1�Vu���xu�բY���Qh�d,��DZ&��Lx�]!�u��[L�N���H&�R<X���4��Y2`a������¦Щ�����ے�$0H� �8�	�����E�T���R�l�\��f�h^V�e/h*�F���ƍR�	��T�a��vhyP���,F��%��#u��z<�rT�Ո9�ǲ�p.X_l�ueB�-������lcc���hi��Nޡx�H�B��6Q*Q%�c>��A����8�F�`�:��i��Gq�j0�ub�
�kk��&a[�i�f�s�,%�����)7����I�����"�Lu�Z�>{~��h�{[�T6�={�PbK�	�,�;�b�e;U�r]ox�#�0��p����B� �<��8]	�͠��@�t���Ս|U�%�29lET|H$�l��"c�m&xT==����I�P%Z�}�G)՝�ը6�8�-Z�@ޚ5bPK�C��V�D��8XOb�|x�����!�4�dP�hX�)�`��fZd�(
��oms�j���CF2k��8X���MIiD4l�д~M7[�5��:A�����"�\�6��b�b�p�G�мyV��Nd1`��$����v���S�}nPh�_�
X�30���oH� �F��PX��,:$#td�E�0J��V�5:��*r�Q60{�^]�MW����\'�D:G֞X5��P���c��%���tH6P�d,��4�I�hW�`v��M:O�ŧQ�\E��n!A�� gO@�g��q�����|jTf���U�V����kd�	�&����Ȃ�S���0�I��������$�4}��Y䲙b��T�i�o�#F�K�A��Z4#�2ӝl,RD�@z����nT���f4��~�Aw$S�		؂��