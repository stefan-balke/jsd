BZh91AY&SY��� N߀Px���������PXoa��� j���!�2h�#������5I�bhh h   @�j�����j{T��4�h���0L@0	�h�h`ba"@����ML��0��z�OSF��B� {�$D	Y.�A�����ė� šPİe5�+���Y
�.�	���tH����I��Ny��=L��o,rm�'߯�j�1WyD��R�m�Ӥ�[��u��^�U�#lr�K.���JB+�h2Y��#'��h����wLH���Q V�����k۾r+��K��$�=��û��;Ų^�-|[���MR$I�A�t�%��r�"�D��^V�+焭4��h�a@y*�^�@�mE��3D)�J�"���9U4h��ŒJ�Д-r����b(ý�W)TCV@�ɑ��evK(�>FC�heg�Ԙ�	-�:����61���6�m%qp���R\z��B�v�
%J$��#c(��(�^��)�(mT���TB�f#��az((F����&4������<�W�6���  ��$r�΃ӄ0�q����OŰ`�p�4�4�Y����U��=��fD�N4��hћEڦ?�I/�8���s���9�w@ľ.�06"�/��d
��Q+I1�Y��h^>���h��3f��@�����|d���f%���&x�I<����_���.��C�Pkd"����Q&P�å4!��L��)T��ypC����J�j��6�}�H=��EƳR��%�����V���r�l$�đ�Q�꯬.׼����IM[�״��)��gf��];C�v�Y��k`@@F�Xhu�y�چ�VM!tWp�w3�G"������Ib[Ҩ��L2`2s5a�g<	�ID%� @H张�;c0$$#�����[na�eI�*��60{�#ս	���%�qD�fGѐ)G�]����dO���ԍ'�C�@ЙN���$�|��&��c'=�Y�ҙ㚼��y˃�^Z!1�� g#$1�G��f�n��k��WI$[�18]"��Rz0�PJ���`b�����H-a��),������R��33��ٛZM#�A��lL �L�ڰ*�"� <8����-w��CH�0hW�v�O�]��BC�6O�