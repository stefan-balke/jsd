BZh91AY&SY��� �߀Px����������P��(���dДԘ$ɑ�C������z��h����ODɢP �@     		
j��6��Sj<��4�A������b�LFCC �#I D��Tl
fJm�zMOP  dlY}B�.���Jw�:�6��0Ш����g�͸.���3&4v5T�`��W�r�âp���ft$�x�R'�W�J�/yT�JD)R�IQm�(ΔL��#�)K�3�=��Xv��DD�GlMt!�|M����Y�s�5��s./w��	de��X�kݐ!�<�/���_�g�M�L�6�wl�6�*h�H׽���"��*oK�E��W�l�ͮ�w4:j����6F���̘�eW*�E㨰��t^`ܾ}y`�����a� �gf����ZP��U\U)���a"�d�䔖�)$x,&1ڡ��Y��{Z�aT��vRY՞�
ɖ`�*�hf���U�w�G�؜��}-��ڳ<@Έ�36�|��Ӡlcc��m�4"�X��T.��9P��犉R�-{�A��*��a���Q�#c���1��;��FF���V*��m(��a���� m�n��7��g�8�'+3m�{B�1ё���i�<
��)�@s}/&vN����GW�$B�wzr�i/��;�m�qZ<�CdG��r��L|Om�N�DW�P�`Td���h �6ۙ�<�㝙��n�q�tL	�ȎOly)��dc%8P�?��Q�`�9P��Y;Y�Y �1�:"�SL�];7�P�2"\�ֹ5t�t�1rL���`ֲ���O��8����N�D6���i]� ��s`,i�4-g���FF�������#���R�ܺ<�Go<}F��l�	��{z��H6!��ۏaX"�6`��G���G��T�B�X�sݸ�W�qφ���3���up#�����uo��u`ir52['z�Jؚ�_{�h�U��´��{�
<<TAb��tHF�d�E�P�3�1�el4\�}d%� M��O���%mǨ��\�S[Q<W-#����fm�TXzy��on�O	l�zpWqԨ�˛��2]\�rTt��ߴ�����id�$�����b���)Ǌ�)K�]��*jM{�ł�7q�Lm�8�Mn9\�~%�=5�\�ZnC���6����тtȠ%!3r%
3��ǳ���-���&b�+L��g��MCl�2m��F���,}=���f-	J}�L���w$S�		>�q@