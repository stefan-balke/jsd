BZh91AY&SY�k�� �߀Px����������P�w]�8�\l̀�P�$Ќ&����OP����h�(� �B"� �      �ȓS$��4�d�=!�z�  h�& �4d40	�10Ui��0�cT����z�MF@�F�2=%�	!�
��T��@����R]t���A+�=�V�4{�S�"�(;�%H6Dl1]�&�z9tt�;�ݢ�:GL�5���`��^2L`�A�@$1K��$�m�R]�6��O����K�X~��eE�\��:.�l �;�QD��Q,h�:<�/Yݮ�"s���c^a��'Ɔl锰�u��z)Z�0cɏ�Xn�ʬ�,e�$��9$ȁ(�`f�
��Y}�6^��B���Ƃ��%7]�GeA�Fb��S	b��"�d�\f-Eʒ��&8���8�D0t
�{9PEA ��K2:�X�"�RMr���A[8��5 B���PD5-E�LB���C�׊��UJ

)j�����m�r	HBZI%�3��\�ߒ7lrɀV}���+
.��
�S2#�E�YRM��`MYY��wSmE�,1�ea!! ����~�Л��o����i]W���l�˚�{~��1� ��>�x��=Z����)9LyO�Υ�������t�E2���Ӕ���,���4���9zO�����R�ڤ�P�h|����Ί������>Z ����7�$�JZl���yz%�F�|0�I����w27�\�wL%M5�})�V�g5�cu5�8��N��E�J�@"u Q��' {���}���f4F]�bP�
O����0-�>q���7��["�P�����_��"�����X�GN��o1�ܕP�h��ʄ-f�I���Mt;��;o��u���y���-�"-]���i���CE���[m����&kv���Cm�w^�e�"��4��ajL�]n��`4.ul�!qU}�U(��=J_�Ľ[KzW&�YXRac�b��B�7�5��B'm���y
�jy�"*��|����u7���
78�+��6&+��Y.�'�i	�(������W��Ń3����F;.	B�q�'�����,���s"ԅ��g4���
ج]8��/Af{�DҎu��hLR�^f��&�r��0�H3K̥�i��W���G����h1����d5�
8eCݖ����E�f��h4KNz��rE8P��k��