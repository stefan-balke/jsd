BZh91AY&SY� �߀Py����������`��� 83�� �SS�j{JyG�zM�ѓjbz44(��C�  � ��L�i�����a�0  �ēJ� @4h4M �2i�# `F&��4� �D�Md4&��M!� ѩ�� O�$ �� �HP }�/�r3�Ђ�
Bh	�!�k��m���+F�`�c��D)6�E�k��t_ӿў4��~��M�kZ|�̇/Tَϫ�@/�4I�#���q|j�y�C;��n��A*�s�݉���P�DU�ќ�!s�a���Śɩp�3f ʝ�SK=�5Ȝ�b���i �[�JQ$+�-�����C��~��٭�����ZDTPQ\��Z
'V9%+� ����D10��w,� T$ f���qRy���xPdS�S�����Z�������BZI�li��mS5 T�Uu�*��q!��)w1`�2,	�'�	r�%U,��v�*L�UIdG�M$�:!b̔,A�;WT�+�-:�C�yd�/�ְD`)t�t�Rmb1MK���K8v�:��Z2._8mK(��2섹#AF*��,Qˀ����L�=����XffQ:-4�hm�dʪՇ����C��'e�	�Ң��҅,���&�Y��=�8Z�Fr�w9���$!!	r�I%B
������ۅo�8�P����p�j�
�������]Dв���IV��#��@J�RE(:h���E���8�z��U2:G�QPQ ��b���P�;��"��=H=���O}1����o7�����(�k���k������ӯ�ӑ�S��q�up��W�G���	��s��Y��>�#%�� ��.=6��{�P�b��$�yg=}+�g��zK�*��#�&���B�3��b�IX��f$�����A�S�I�@�k��`0c��i=LōA����Ֆ[ڠ�Q�ѽ1	��!�Yb��*�L�;��gϨ�^�����m�1	Ƃ���+�?p���CA��LP%��o�L'��i�Ɔ,dל�7؎���a�1"!�7���#����W0`����A�ya�.��V�#u�,ZD�|���=�oۭY��ӱ!ߨ�G�C�9@j�Ztr�9�A���\�'3 �75|�q1	fG�L��%��U#�*��]��e�]��`��P��!"&Ȁ����bƚ��7�fr�#˷�`zm3��� uq�H�mX`n�1􆡡2�NFఐ$e#��h�a���HE�1=�����y�Aht
�}B��Q�聛����lK�KNbREG�`�����ͻ�ha�e$XH�'P�7n^%S,� �4�P)5��p�d��Ae���%�<���r�[H�����`����AkA��͙J�_$@͸�>r6�͊�Y��fA�`в�d��ܑN$F�1�