BZh91AY&SY�in� �߀Px����������P���i�iMXI%1O�=�<��"dhhڀ�  ����4�P�b0� �`"�AM�hh4�i�h ��0L@0	�h�h`ba"@��6��ɓS�H4 ���Ad�}���E� ����R�0hT0V�N�s����l2S,�;����Z /}<���e�Ɵ���pj��[�DDV N�P<Y�-D�JJ��Dc�t��g��{ur���������8�n��\eL��G�>rE��5I��7�94C����u�$�o�d�
�e��������~�����<�[�i��ɨ�&Z^Bܷ��^v�ENrP�C4�����(� 6�8"0:����L�-�cܖ�xA�44q��2�3�Mf�c�vUjOy��I��B�6����}Z P���P����k����,�Gh�UÙ=g2"r,�d�6@��f�T:Y�J)�Ȣ
͒�p�y�u���2aZ�@bH(!��Ɗ�2�cn>	y��spn�j�U�Y�3�M�C����61�-��CHP��� �и��B��8h�(�׻p.�1l-9����!yV$r&$#iҁn�H#}�Z�eD-�e�B��&a�-<�.\m.�|�����v����$.�?}Z��\K4Uߢ���y���0�1��̱T�]�Lҟ�sv�;A�ɝL������5�6Z�xcv`�O�B� pP7��vj�X9��_�DWvW����,�iq�Yѩ�'ʡT������4C1>u��A�]ڒxP%Z�}5�捧Vm��Pb�DP��,��D.	�dР���.�P��=RЇ>74���@�cll`�`P��
����{��5�)���O��i��PB�Ɔ,d�Y$edts���<�H���dIhU���#W�u�������ߣ��S9X��Y�l'8�`L52I%�!����� �(���=�4z�����m1�K�p
�EK�kCs�oI$�@;{j��A����K�\2
��b��ju()4T<KQ6Dg߁�	�M�a�0��"��x���ﱤ�|(�}po�3����1�#Be}G��,I!> j���N��4L�>z�b��/�MB�!Q�聜� ��|�JA�rQ�|��p���ka�f6-"��Rw��(!T�&���ph4q��ȠsT��Xh�7zժ�P��"~&�����k7M.2p.�Q"�+1Qj� ߶�ߝ��nT���� �`d)f�.�p�!N��