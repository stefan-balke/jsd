BZh91AY&SY9�� �߀Py����������P����w�P��GTr
<%�MOAOD��h��h@i�T���DPɑ���`&�� ��!OS!�#CM4�z�   )CSHzM���     i��$I4�FD�L��?T���)��@d@iSB,g��*$�JT	�#�y�_���I�2���[6����D�0�Z��5�R -}9�0��O��Y����vd^1��EF�j}`4-K����UBJ��;9>�!O�������ƮNH���b��.Oi��*O[�D`��ҵ;�T*��.[��ZB��>�@߮vR�F6^D'�Ȓ�CiaˍɈTPQg��AΡZ�P����]��Fg<T�E*%)$4��S��9.*�^mY}��B#[4:v8 ���rMXk�@q�#��P��Za�y2Q��<�p���ĥ�f��\�3QZ�s6,�����L�$v��X�`+=m�
F
���F�J��ҵǵհ����(�c|�P��mi�E��*x��i�(�N��ϵ�+d;	�z�\l�Y��Y�[U"��nN����7���hh!�r���B��G*	�r�*Q%����T�6�UM�UX�1��F� �PeGTKĎ&\j�*Ah����k�i܃Q%Ҳ�W�4�1��]%��%g��5��yKo�@>�7�Q�T|Hi��>��>Fv��mRv�v�#��եB!�u�q�J��n�^P�r��u�����Ь�F�� ��!�eUc�Z��L���h�Q�Afj��I��.�a�A%����h+?mF�A�,�I<&��-�(c�鬼�Pv2���K6�	��1������uf���8�B������M �Q3�`8"�\�LD�d�h��o���g� �\x�{ eK�$s;lDz+��� �4*���lq{ ��	��20����|�:�zL�\-вhP�_�Ax�W]i�{�łƸB��_G���{�Ʌ�0��XJ�4�
Ɇ�Ъ��)ՅN�I �� Q�ؠ�w�âB4/a.�p�+o��Y[⦌�b!K2@�w� �ڄ�.+��pA03B�����Xw-(�8yA��uA��>���d4&�x��BH�qM�i=;@T
�Tx�(wK��ΰ�@V6��3<�Hc���I�Xn�Ɍٷ<\"�C;�bgJ(�x�<��.�ΆB3a��F�����:�-� ��s�"�0�Q
�Q�Υ��1����4���3`Z�d
E��hXIo���׸ܧJY�3�j!��B�9y���"�(H��׀