BZh91AY&SY���� &߀Px���������P� �0*� 	H���z��7�)��OHѓ!� `LM&L�LM2100		"M �d 4  �A�ɓ&F�L�LD�FS�z �!<����=@� ��zG��Y ���t��$A��������0ШhV!M~��]��aA�d�cMړm �@e|w�8a�~<�g��mgT�'O�u���(����e�1��c`r��7�pg��S,aC�s�ZArw�3I�'1h�O	�z���M ,�g1�P��g�hd|�QW��Xe(A4����!��ʴeyK��{���գ�)c�/^���++p�����lY并0Q�Pt����G�$�cc�fQ2����Lѝ��� ��˔R�����]wehDC&�.2�Q�ښ�9/a_"���h��ĚV��UV�E��6��lcv��m
=��_ �\<r�Bw�
%J$�c!��rUe%��#V�TfE��.r�v�a�P4�gE�`���1�m$�M�}3�<cF�6@�h:d<vx�]�Ab�挶aɡ�O��*�k���۾tj��M�)\�AJ/��{�G�[ ��}�^�<�)�p��4��`����s�3]�S d.frBƠy�l^�2ͩ/[�Px��F,��
	��W���6������de��N��[2`U��Y��nnƠ��E	q�65A2���Rhn0jإaJ�#ɛ��t"$3Ӊ��[̄�M�J�F�EZ�[T�G�qp'���T����""���:��5��&}d�3�	�1�[�ș$#F`���$�6��DU��(�^���Zמ�Hh�`�,k�G���{��g�Zp�	lEF����b���9F��#v*H,A�Ą�i{It���Xa���b�J"M�Q6DX]��w�By�i�L`|�$Hb=���_��ļ �k�>��r���a�2���hXI	��z7�3v'-@�
���*�ð�2�d�P�xPm���ɪđ1Ţ�Tl*3>��
���-W�,�a:�Ԟ[v�R�&@�:@\55**K.BAe���0��)�i�=W�ZL"�����R,3�J��$A�\�����jZJ���3Y��F
�yi���"�(HB�]R�