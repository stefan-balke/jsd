BZh91AY&SYKlf> �߀Px���������P��r��L�,%e6���j#j4��C ���#�@       BA'��L��4  0��A�ɓ&F�L�LRHj&�OS�F����OF��Hh  h��9X��҉,��B�W�������1a�@i�&S^���n�d�j4�dCG��m�Y�5}�'_W�W���=��G�S�ΧZo��D����^'�xZ����fY�m�gnS�pJH��9{G�����,`fJ8�כjCd�is����Q�[��o\�����N��%Σb�2]�X�=W&�0���Σ�pa@EEr��|�BD�A.ŖƵJT���wuLG�U� �K��Oy�&KBGzі�4M3C1_T#�՘z��xD�#B}̉(�Z�1�>4�-�n+FE{43=�K
��L�zJ1+T,�"�˅����3�aӵT�c+H��5Zf��3�"��*�F��U
h`H"��9��xA$LLL�L`%0����l<����a��<�&�&��[%�7nL����u�lc|m��!B����C�Iz{H� 'y�T�K�X��V*S��֫�L��YRv�{oK9"Y0^���<���ZҊ
�廞 ��bM�f�W�C3��Q��K�����3��N�Z!�0a$�Wz�!�����-�����=�������U� ֵ�"Qj,��^EJKM ��Ę���5�4�	_�B�Õ�]�S�����O�)3��4o�x�b���x��n�%JtP�?�0�J�-L��],��g̒|n�gM�66iw����P�"�v�<\.#���3�E����`��vcr��2pZ�`�m��@�"���*���a[�ns��6̒��z�����۶QP�X�'k��8�_�Ӌ?3%��D����T�*��N�3,%�������9\'Z��bŹ���^[����"�\�YHg}�7c�*:��MQ�F�a�[C�``q,�s#v�j�K ������|K�}�E�P�3�M
��Ū.x/"x0ʘX�3�w�ĭ�b���Y�����
G�G��{y]�޿fw3.�q6*&k>N�I��'C�
QN��)��o��dL^;g#C����M,��˪��
p�
R�h�V扯��S�i{E�5n0hcrʞ�s@�mD!!��o�QI�깩�Р�F��p�]/�W����s�)'г���rP̘43ƚ�����}�u窦��:7�R�1�APIg1���w$S�	��c�