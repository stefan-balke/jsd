BZh91AY&SY�}�� �߀Py����������`�C ��AR
��FI�OBd�5�zjze��M= =A��JS��&��     2d�L&F@��M#4i��)G���#&L& �4aLFL`�&M4�dd�т0�F� H� �������h�d�4d� ��4BI�H���T������M(�hR��@d��?�6�]��\e�@����rD �_W�p����x���^��1�Osn��A���$�ӻ�r��)��|��d����T8�6Wz� ��⮌fe���fԗ5��+�0��ї4�M�Lf&
��NO���vƅ�\��:l�� �=s�j)B��7�6�JC�H6�}�4��C��U�: &�$��������:���hB{أw�q�z�L� �&8}��,:��r��[��L����v�v&12���V�U�4^�}��L%#WM%�4�A�I1m1b��L�5Md��#F7�}l01L���n�<+�%%���4�`H3Ô v�.�$�Q3�H��=RSY)��(L|��ZpKp��ť��N��8g"b��ӂΒ[|�P�&p`1�EԦ�Jk&��1"SU��b�=^䛨.�T�H7x�By�e�cc�D�ڙ��ٹ	9�/sߊ��k7�EWO��^r�ֹ�M�bYV��ꖉ�`���5��"����Oj���U6��ʖ�&ܭ���d�E����h��C�����!��"������X+Mޠ�����*j�S`U^�v�/�𳂴��C��61���m������|��E��!��)�v�B��Q�`�BE�!�0�ɑd�'q��9L`w%�"E��.��� �rM�Ri���S(5I��@ �䐐as�����/����ǫwM:q��A������d+u��=�}v�����󂀦!Dn8�� �1xv�ձ��;!ϕ��\: �o�Ǵ����= sP%��mKW ���k`�`� pD<�'=#���#h�HPbD���\��b�d��%T�=@%��PI�O�Y&o`s/����d3��X=��Ay�Вz�ka���M�x4�����jVB"��)��RU oh7���<�5�W���\ȟ[<xQ{���K�6��m��C��N<�p��n�"|�� XNV�'	:����8�:*mc(��9�'M���y$�m�ѢW�\��z���=R<�Q�7?�lu�ZY��Z��8��7��k&�_�(��� 9|@%��; h�W�~W0�N���`J� ���@����-�U�R@d@q֠D�o@rD��U"��R��^�EK�X=%�%d@F{� ב	����f �1��2G-�3d�"�J�>���BU��7�-	�x�À\�	dG5$�q<� �Q ��ֱ.t�F�,8X1�+�T�pc$c(�gc���(���Ѝ��a��k���8d��y.R�E/�ʀ������l4�C@�
Z�X9�c���i���F2( `�)F^�.VH��_Q��d#����C&�rA&�`F��D�6�{7ٲ�2��6�,,�с���O�rE8P��}��