BZh91AY&SYW�0� _�Py����������P8y%C0Ѡ 	SR�=)��L4!����Ɓ1��L�i�����a�0  �5=�4h�z�C�h2h  =542i�# `F&��4� �D�dC�Dhڍ4 hɴ�H�愈HR�"_?�rt��4)*d�����5�B�Ь2� h�2���w�l�N�s��>��v}��d��{�U����
gTQэ��en>�A����C}��TeK-5��*��,�䌴+M����{+܃Z��w� V��P@���=�c4�7>�e'���P&�1�}�&��a�s����zyfY��ɓb��AsʁEW!�������H��ch��a}5U���G{�i��m1�Y&[��f铔(�1���tJ%�M�Q�]��z�ٔ��(1�C��d���
����B��m-�j���H!X]�c�t�4��lc{M��CB�:��	'&	C�q�DP�X����X�d�)E%�Ô��@�V����L䂖�BA�5���M	�b�FR���>�A����R� �yS�����"���Wi�P�j��
�B(�8�qO ��b!�q$}�Ӝ�.�NwF�j�l���{�WyF�����~�׻��J�0vM�����OO"��ӂK��^�_$kf�ƁD���޿�&1�f�¡��d���'�U��S1�Ѱ��`X�FB"�s��Pʥ��ibPNb5�Ua
U#�9W8���ݰ!�8̡�hX��@��pk-���%�z����9�.\�nc	��H�b<�:������h�SBb^ea�V��d&!�[/��n,`*�+SP���1�ֹ�h�-K*B����; h�S�}NPh0�X���,S��V�Sx�HW��Y� �������D��*�B��ju()4T=%�Q=��F:k;tB{��I�Ldb"�D$|��C��#z��"@r�-�9�Ik8y�>�hL��wB�HX��� cG���4L���I�\A]ơv��6�0��d�5��'$P}D����i�fB�"���H��BjN���R��fbb@��A@�SYu��m:[�������F��NƑ�����Ѥ���s�KB�DH�ޯ*,��<�w[^�R�.���6�y�@B;�f���)��Q��