BZh91AY&SY(�F �_�Px���������Px�Ց�q�Zְ�D�i�=�����!ԟ�4h�z�S�T�I��O)�� 44   �I�A��2i��4  S��& �4d40	�10�!2i=)�e6�2  h �}Q ��, ��~�
m�)�m@寴���F����r0�H/�}���ո�һ7��#ﰝ6-���u����]�'#<U�0`�bk΅2��'yH�ӑ2O���� �焄#i�A����N�i�_޷5�:��HLy�=q%��J9#�\͆�
Rt"�2�8ʺW�"cCݐ�l$O!�s��È�u�a�PE�-�\��HAhǂ�C�vy/�I�($�E"�	�Mb5�B$VVZ�VJ��[�{,�wѓ��c$f���{���A�w����9ya�)TWj�#��L�;�08������1�40��Ol0�NeO������K�>�_<;L,�l��z��^.�Y�����19���'�9���R�u�|"�>����q���콺�~H=���.�Z��H�Gr�.�����p
�N�q�f�J�mqm;����N�`�o9V�`�1�@� E�8����d=--&� �t���#e��c޽��`�h8gT��s���5�6k`�jSMd�\��:��*2eDr���(Z���ͦ*㠗�W�~u��X�JF$��-����3�7�S#Dժ�)���0P��W�JD2k�f&(�b��N+փ4�TX�9����1�h�-.b	�Pt�;Bf҇7<5����J��u6���!����|�B�9s���s*uG�,�Jn��:��j�J��]P=s�� ���^��C��n�i'�NǏS�)��>��A&�?^���W�a̛CY�Aq4?���&�������(f�L)R���	{�T���kZi�,�ED�C���S���F��F3;�V�1dR��1�E>WCc��]�"
��@��PNx�GP���ײ�]\�1UWg�t�(c�����)�F8
0