BZh91AY&SY#��� �_�Px���������P��8h� J�=LL�M��& @4��� JFS�Ti��C!�  !"	���4�� � 9�#� �&���0F&$22	����I��Ph S���SB�'������P� {w{�F��q��(S_���8m�1��a���j�1�3|[�W{���IOap�4�#�G�E��uYZ�����'�*q�>v��s�d�;l�eFXL�s�/����f��X�+�Յ
��3,�+�0IW-��X(�v��u~>4ѐ�o�;�}�����dZ2	��Ih�MH���ʕx���ay����i�����6f:�b>bd���eD-L�5c���#� �5GTbI W�"��G(��Ԑ�E�(�EP�(��@�)��_j);��aIC^Qd�j�2^+�������m"��;a᤹:�r�R�z�R�%�{�,��S�ǃ�n��62�8�QP3�Ψ(F�q-��Z4�==)��;2��-�]�H�((?���d��B��hrTv�z}�Y�o5A�2�����F���&�:Y��%p�L��$}���_b�����[��A 0�e�w/�)�pL�H+0<W���μ�\[�%�^`�Dgf��@����z�&1���P;�2<K9$�j�[.2[b41/*�Y�.��kTC(�sB��D�����*���y:չ��d���+���3�橜	m��(!�[�Be��D,p��-�0b;$B�$�H�8u����L�5CI��@��4lC(�(�	�����(	ݙjb�����P^<��ylֆ���4�`��Gh%x�a��q��XKhT``L31Nfp�7<gy9`Q� @H�ΠD�d�K��x
�s��Π̇k&�h�XTM�My��OU4�����ǻ0�G���CY� =���6��g=�GpXI!�!ut��# �&z`�,8KC�V��B��s@�ۆHc"Cd\���aA�5l�*�I^/06["�u	�;��PEK�2!�̫(^55�Է%�����%�Q$�e�ɤbc���s4�^]f���̉�e�E�IA�l��[^F�K-���i4,�Om���ܑN$��@