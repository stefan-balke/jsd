BZh91AY&SY�J� �_�Px���������P�v�A��� �p�BR{JlPi�4� �Q�� ��i�Jm@ d     		iI�S��=�zM� =@ �`LM&L�LM2100I"e0M6�ML#S4�=M� �&'�ҾH��hF1%������U�r;C�r��)uO��_UV>�B��3,"�q������Gw>�W����ĻK���\m��<���i��d���E�����C4�ufy1��s.ްu����6�4`fIJEr�w�IQ`A�!
H�!L#���h�
���,k��]Y��b`��ԍ�{X����W��{؝hR��+>^��G�ѢpgM�z.�f^�9�R���iW���]��؆M�yV��@|�)ɛ�Oꃽ4ޝz�5^��P���ζ5X�g+|�Uhse��\��N]��{V�wT�}˲���V�B��02L����$��ֶ�\e�d�f�D�H�a�J5)�B�(�&44`��8�P�c�:��<Ncc���CH!w�;���)/�Aʅ w���]��ԑ�H�D��	|Щ��N4����2�7�P�(��aׂ����{����e���K%��7n��_�ux�Gfq�s8|�W�N���S�W���1o�$R*�Oo�e���}�թ�t�=�䨳����?_F���?�{�qy���,q�^Z�mӵ/;�Z�����g�Ly��<�LUPw��)���3%7��az�JZ�����HC�g�I?%±���X6h=#��82�;r�ڜ�gt�=4�̀C�E��K�*�ުt�*�||lZ�~�"��lfs�ba�W�q��?*r8�9'ɂ^b������6ݲ�C��qt�<#�Ǉq���z̰���_*��{4�k��K��4}5�n5s�����C>��"ŋi��0�ߺ*5Mu$�pއc�Tt0�W���1��l�b��(q�5�)}���n��S�� ��@���A �bBB1a.�p�+�FI,`�#�����V��z9�V\�P�x��S[�֒�#�w~'ݭ������79��8��+�6�%3u:�#��5����S��zн�gb�y\GRy3��R�B���(f�Eʵ�Ӿ�����FN���-���M�����P��:@p5и�����ɿ(6�h<֡t8T��F�TB�岂�DT8�C�( 4��h`��E��,{�i����fǋ���C%;
�O�w$S�	��!�