BZh91AY&SY$ʴI �߀Px����������P�wMہع S  �E6���L�OQ��M�h�@�4�0)H� ��  �  	L�4S�҇�$��z� h���b�LFCC �#	��#И�Sɨ�56�jmM 4�������B($�����0��
I���&���m��Ѓ@Я��r��hn.�d�6��m۫b�Ե�]ص�c����!������BY����ZT�*�MF��uZ�$)X��g;�Z����
0sAW1�̡hp��5ٔ�W�C����t��q��QV�|P���v�1"�_�V�t㲕� ����L�Xu(q�`�K�|�}&^�؜~1�y+�C1q�1ɜVs�J�R�}�@�Py�D"�U���:`���"_R;3\����h�b ��Fm4�hP��!G�Q��*j�+��fU4��W��YK���DӺ���4��J��k��T��sD��dB�b$+�fh+��7i�����H\TC1x�V�XNe�0v���7�lcx��mc8�׸:�F�p�s$����r�n��KQBPT%�7�%6�n�hE�J�%#����T�CT��`e^I	k��Y 6 خ���ߗ�=�״��n�q(a���_?y諴h�Vt:�����ǟO�H[	,�_5�r=H����6&�j;b��L����l�3`�5ۯ^��yG�;[�4��A�^u>���1P6!��}&�u�3^�R,�c�$�$d�g�ҡT���E�MC3�P��dv��$�4	V�4Pԇk����5l�E{���� F��ohPK�C��V�zIw3���gנ��]�$�bN59s���A�ј��/��T�Y�ύ5OR�i#�衭�&�I#����+�{�gD4_)�f���Ql*k���������M)B"�ʔ*Xy6R��,�o�YRԑ����9Jt��:��4��*$��s2
�s�oD@pl��V�
FƠ=��@�A�&�防�n��X�P\<%�!�"0۩��O:q��I��L�im�ݤ�`��/�f��Fő����Ƅ�9�ÀXH�@�����ױ$dg�KAa�t��@sG=�v���t@��Hcc�Q����#yQ����*�+po���a:���p*�*\H�"fx�
X^In(X�.��Am���J��3V a2dei�S�iy���LGq'9��4��a�\U2D��w�^��6�Yf�G�̆��`Я�o�.�p� I�h�