BZh91AY&SYŨ{� �߀Py����������P��y��u�9h$��S�m4�hS�4@ �*h�I�$ 2  �  !)��&��2d�M�  F�ISP0 �i�   � ��24��Sjz��ji�� �24yH#���l@��'@!��F	P����:�D �mI�`$�M��K� �`�b�A��R�H�1�3m���\�0\{`a�:D��XaX�!�/�-R�7��Xo��L(i�$�wxޓ�E�l���6��o4ʰX9��Ȭ�Y!��yd_�\jZ���V|������������� ˮ���_Pj�Y#c�R,��Ag8��d�0�귈3rI5��K�7>U�U�ُ��!��<�����!��lK-g�L#�wC��YMd0Q Mk{�Cyk����dD�$Q�`Q\[
�<�MU[E�
$�e齑��	�م/&�H�:�U������h�	!�B ����F�M�T���$�YYQ�a_/}�Ar��c��m�6���8�j�KĨK-�'B�vS��QQ%��j�mT��U60��E�%�Qْ�P�2�	p4R�@΂^�Eѽ��lCci�ik�i����͕�L���ôqs%�^=^�Ae8,�՝T��K2�!�KA,�x��ǅ��(�h����&�RFj�:Ǥ����`A�)m�US(���X���$�LA �Ց���4+��0=�����}�~�в>�|(8��P3,�xo�p
(3(U}}�H��0|�� F��}M�CB�;7�ȋ�#8$����f��U`���r�+RC�
+^*�9Vd7!���~�l����0�Iȩ�0�[�F�R��ϫ�o0rJ����п��\��  ^�d��	�ףi�})4(k
1��L�؈	�ꐙ.2"�2�K�s^�[�4O1H��9�,�A-��0l#}�Y��: �78������HN��itNA�P�vX��.%��@V� /(�o�9bQ@�I	����T�0$$"`z�a+iy�1a����ܢI��zK J�JA-�<�� �j�/q��˸�'���������'	W@�d����Cl�� 0��Eй5c�V�X!v����(�<2uô�t�.Щ���"	�@�$�"\�����\��6��̒�GXbiy�(�(�5k�T[��څ	��b��d�AP�S�K܅�+7��&�	��?C?4��i��,!�z�L�T�f\���4$i�A�i�!=�BV�~�d@9���l+���"�(Hb�=�