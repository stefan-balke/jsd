BZh91AY&SY���� �߀Px����������`��)�s����~��C�� ��M@    �*L&��Ѧ� Ѧ �0L@0	�h�h`ba)�����z@��D   9�#� �&���0F&$
h�)�S�l�6�&�M��3SQ0� ����$�>���9��U�HL4�d��I����4�hV,�;Z��D	+Dϫ�{�黭YY5Tp��aV����v�i�:e?��拡�VwBw���6稑*��;:�����qd�R$�詿Η	�Fsy."��Qoi�HН�:�$Re5��U���)Ôv��lw��! �����hH���&5
b�,hKCm��V�s~-�O%�d@IB�^��6��)���8'lƂ�_m��X��)q�1J�O�q$2>"�4�|��i$��RS�5;<؛a�^u6Ƃ
�9PT��A��I(j�9��eQ����]Z�ќލ��b��&�a��Ƭc&҅�,�"�|�	����,���eJ,UHq!�$��yķh�ڬ(�%Q�Ax�7��*�bb�	�j$X`�Uy�|�	��akgt��+R�U)���( t/���Ĝ�D�2���Zd��]=2��x7Z%3b��f�C5!��$��I�j$�A���.`���N����%�$�P �c8�pq�#oӖL ���r�n�uIؑ�S��11"�H����tM����It��I�2�w"��32����@�p�V����������8C,-V�� �o�â�v `fN
]����Ǳ���� .PHvܠ�d�K����DD� ��"9�$s�o?CH�ځ���!��������x|��q��H�BQ٨�Q��h���� �����xˊKʑ@Aܐ4`̏
g��	��m>�w��A�h�I<. �Nֺ��X0i٠657f���DP�Y�D(�fњbC%�!�Zb��It�������9��b����m���q��a�,��A�fA�h1TJ��>��U�x��=471�ZO��9�#���A��L�o�5�h[�i��U�1SW�3j�� Ժ�m�ܐ�z�������>jָp�Z����@wv`:
u��r��@���Yb8�P`k&��b����H@9�P"A2[�R64@{G%b
�B�Dt˱*R)b��EC�Y"l��o�#Ͻ	�Ā�3H��^$@�<}7���nZ� u��ddp�F��9����2�����(� �����>����#��$-*�ׅFӢg�"��q�B&=bXp��ݿ=b�"�zR03���MIݧ�Q *i�E��j&���.� ����n��0FS�
1�)yZF>/~&M&�wq�n��,e6i* �H��P�:]�I���ᘍуB�挅ܑN$-+�� 