BZh91AY&SY�|�� �߀Py����������P�׮�u4hր	%�jx#L�#@h �L�������"*0       BDF�������44�i�  �@dɦ�L����0Fh� 	L��JlM���F��4 ��h,��Đ�BF"ɤ*=����p�A�B�Ь$E
k�_�����8бLńM1EQH�d﷬�٧�jҙ��Q�������(A��x530��W�QMΘۮ}��l�6��b�u\��l��z08Aaq�t�^A�w��$H0y뫜�H0Y<�퐄�e���H!�n���M�C��T��hhrX���B�00����B�&~5&��ח+Y�ծ=��)v��[k���kj3wa���+���݆��1�G��D2]H��h�T���}]�"
�CAb:<�U`w�������� Q!�B�"he�q-%X%P( �(.'CF�+ ftP
���)D��]�]�8$�tR�@���;;	T��
�#��� /�]�\W��7�^&%��2��n���k�����m$BW/�Z	�P���Z�ݲP�f#e�3V$&PƩ�UT�M��2�G,5j���-�#[��!�Qah�f��z�`�Cfh�'8j���O�S��T8|�Φ���W����a%�6ɟ3���E���4�4�
Ņ��'�f�Y(IC`�z�ެ?^�9��ď�!Ay����n��h��j�N�ui��K�X �$`E�)4X�	AŁ%�"la�yT=~�yoD�Ɓ*�ڗT�91m=K��s!C�T����D�Q5��![0k)|"�	��Cpg7"���Di6:���^�� ����Jb��T�S�|�����PH��Ԗ�5�MlQ���3�$AtF!Έ[�3����� 1����n[ B�"��T2O�}����{+Z��41kX�o#�������}�P�����A���`Ҝ̂����*=dЂ� ��Gױ@��XtHF���H�d�:f�5	��_�E�� �l�Î���	�M�G#�S�J�R#WF8C,D�*T<�C�&��WQh��A��Be���y��I"�:��M�k:p,	�g�J��a�Z��J��FӢi��fh�D�^JH��\cB�3�!V[�K#K$XH��B�ں�	5Hd̆``@����Kn��Y`��n���1��F^*�F_�ᑛI��i�o��"�5��X�i�٥�y�R�-���"n4)`[���"�(Hq�J� 