BZh91AY&SY̺)� M߀Py���������PX�3p�� %
jOԞS�H4?T=A��M ���h���Q�    BDS�=F�d�F�����H��2b10d�2 h�00	#�Ҟ��G��ꦘ�)� �'��H��"���P@�k������A�B��XI��I���$5X�hX�b�GUDd��d�٣sgt��{��NPqV�����~V۞�V�`�f)���rT���w6~E�q�F�fPP��k����_Dw������������[�! VX�b�)��E����@�R)����q0�cm1٫ݾ�b2[�M4����:�j�QO9N� S49���0�(У6r��)��fXM!�0L�K�b�q�/�9}wY�, �_b���C�TC���E��t�]��u$�v�mb�þ�����_��i*���,��$J�&�D�F'Wc���U��g���A)���8���7���hi(C��/�ZKN��RN�R�/X����`�c�l�.5Q1�B�!Q�$p2���-�#]���hmfk^j�_܍c�b=X F��3c�垛�:�RQj`��Gx\�!Nɣ��L����Ŗ�j�V^�2����z�%D�\`׵b����8�v�&pd
��A�10b$@�@4'��J��2���>uD�	x#c7�&q`o^��I��3"a������'|�4�bY�F;[N�EZ�� ����mM&L3g�4!��H��RU#�Εև��1Sn���'��{��L� �[��a���#����<qL�8�DWR(�Dt�O`Y�D����HY=2�Moԏ����@f�9�ĳv��\�o`@ ּ7���)�|P�z��,���n����:���e0��Lp*K1T``H/`JF�`V-�F$����J��|"�!!]"�E#xE�2Q,:b��P���������D�� ���F#�<e�;m�F' �>���\V�I�Ƅ�vNaR)+�|�`&��cs0ӈ��D�xlW:����Vr�k	��$�ȉ h�HE.KWfPf[�T�)pgp`gX�%@����DĨ]&��5Aa���a�F���q�EQ��>�F/���A�@��d�7%��q@1�$D���Sk�8���ݘ�C�m�O�rE8P�̺)�