BZh91AY&SY+�� �_�Px���������`�z��.tw�� j��4i�## C&&�4 ���ST� 6�     �JF���i�6��L@4�h4212����� �4 � 4@`�1 �&	�!��L���M4��f�ɵ4�Hڌji��hSM$Đ�� ( ˿�;�"�A���U�U��-��}����B�4+,a95)ȀJȀ����n����B�:<-�����1k[��u�]�[�iv�O���*�M��:쪫�6����3�RIgR]���F_�O�- i���$
*0�F��4����5ҳư�!C[q���@�ǩ� E��'4�����p�`�	����m�n!T���'��P8�CL�������J���`�C��P�i
�Yw`��d ôw�O����H�?`��P(�ʓ�*����h4U���|~#���(��B1�����z�&ѩ�ѱK�L�ؔQ+���@��
VH�/2�'Q�K8 �jy�GeF(�b��&� `|K�t!C���ʈ >Ud6@��FGz�p��a�wv �5�J&0Hrn٨d8��.]kAl�7L�CF��Ի٣&(U
9ȘY�aPF\U�[N�����mZJ7F1I���"�0�vٔ>�P��Ф�`��T8�\P
(iPlX�Ӏ�
"����ДQw;'K��������)ݲ\�Le���p���t8���02"��8"ʍ3)S3j!� ��B�L	wm�CYa`�ks�[�4-n5�5����aZE�g]s v 	��z�!`"a���G t_Fz�_d	��>�a*(�2����vەP��
"�)3����ťR� �P��{C>zp9._�}c��a�G���뼉��W�*h2Xd@���x�IW�����KA0A�@�b�c鼨TL���`M��L�dP;��A�Yؒz��l�i���ë^��
��.7FmQ$�$�l�&�3�D�����*��%�g����gA������hC�e}�`W��=�6���1@Pd���|k�)�@�yD�Q$p�8�k�弙K��CE��O�\�0`�{	��x��b�v��d�K�-�/^CH�ֵ�߹�HYWzz�@|��P.:C	f%Q��0�T NF��7<g(��Z�0t�5
0s�`����u��E
��91��-�T�!���*���"/߬ٚ�O��:�pT�A���kLb<g���ff! t�q���C09H~p�4&W��9��B� �I��/�́������Xue��+x�/
�4��d�0�M�"c����ʌ˛="�"�w�gd�	�&��]��T�C��xi��t-�i ������+���	Z�ܧɤc��bii4q���406��XmW �H�~p,�����[�e�$ �`Хy�m?�w$S�	R�: