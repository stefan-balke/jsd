BZh91AY&SYV�D �_�Px����������P�r��i� 	$$j?F���h�A�  4�a �       S�HM
z@�єښSA�@d  0`��`ѐ��&��D�	�@L�m(�I�<�� 4)�=&bi	�I
�,� @���1���*Ф�JbC$��&�����B�L�`��40A��b�4:tph��v�l��k�j❍���4�O��tku��.H
	eoV��"�n�;�82�ov��͍�Xe��ㄝ�)M$�ÇH���V�lH+W-����au(�+�!�i�fo�!׿���2;�캄�G6_T��;�f���ݪ��3��MRHq4H�
U`�&!=�K�#p����J`�.��Ug1(��iR� ���
'g�M�I�+
�a ��,D@���E��Y[lz���%�XF��"ڗ&XBʡ��Y�� ��"�B�IŅbH�`8*)s)�)r�ai�ghS)P�@��X�TN�p͗��{�@�/0o �/{p�1�\�{�DQB��1I'%����7m%���n�J&���F\^M"Ւmj(�Q-3�M`��TM�U"�UDԡ�T�4[%Eƣ3� ff2"��ٿr;��X�m�?wD0���e��Т|��_	ߓ�4�O�t���9��n�J�(�{��[f{��i�6N��Ů7�F@�0^°�:C��!��;ha#��� ��n,ꐨ�Ð8e�!=e�1=$� ���#C6�
$��k��&�2��=l>�Aq}ROEU���W05Z�Ś�[!C�	pj�2�8&�2\�5�R��X�d�~h���F;dXUUw��V����u��@�0�-E�1@P�a�߅4�J�bGGE�d��I�G��!�y"��U
��+���� `���~�vhTLH�~+[A �A�~�굫�%�bδRR�$x}h�:�����y���*���s2
�s�7�$ �@�	�( ���94��J�Vg!t�ju()4T.,�M��d=ې���8�`2�(P4�.����9�x� 9��m9hdp�����2���I�	4``�s�p��P	��+�O��^�_���p��t@�^�c^�b1�2KO�*3v�ga�9p-�X�BjN�6�*a""�%C0ԅ6��K,/��.�`u79h�%T��B�7�R�cH��z�6�����I�/h6�"�ՁT$�7��w�my���߫2c��%����)��Z �