BZh91AY&SYȪ�� ߀Px���������Pr%0֩�40�DjzFG��ɣFMh��4 4`LM&L�LM2100		O!	�M���L�  4�A�ɓ&F�L�LE456�5ޓC)�4?T��OI��yLI<�$$Q Y����{�=#b>�AV�1���_0>P���B��0���j���0�2{xή��M�I�1�C
�Q>�+�lׂ��/�L���ض��xA��ys,�&Xe��#��N�)�-S$i�M�r��C���b�q �-��D�S��w-�$EҔ��Q��P8cm1�/Ӏq�����9io��	)���Z�uʾ�m�3c�zhէN�4�\��'�u�3`]�bx�T�Ҝ%�J*:�	�"�*V��i� f��,0��oKXe��eE���0+E7z�R��b�[-������<�.�.cX���7�m���!�h��%��#�
C���*Q$���`�!f:#XH�$l�M7xZ�;,����B�U��C�`�*���.��5v�fw��}k5��2g	Ɔi�y{B��'�n�!ծ��c�	DB�7��	R���7!��������i����Ę���51.�b;�H$���M�lhT�2I������Ԋ���f���TGh�$lf��@�����|��2(z�"GyobI�N���֝��L�R2d�B}%�TC(鋙�C`�Y��1�lxJ�g'A����do�:Ԅ4��)��,�1�����^r*	�����XACB���j܇��ӉB{l�������]�V��Aă�����|#�BN�QXM�
��s��v�EBu�����#�Y�G���~��*��5��\F�X`b@kb�.
ɸ�'-d XH	͛���|%�	��'�F�[Pe� �$I���*
P�خ��O*[�n��)A����I���\(̓4��gط�K�~��hL���HP�����z�DbDX��'��80h��P�N��YDX/)�-S��f\��*���Z��2�T!Mߣ����&H�)+H`5$�t�����4zJOQ��:��b�ʝM#_�ݬ�i4�ĎA{j&X��TX�7� ���ׁ�R�,�h24i�o��]��BC"��(