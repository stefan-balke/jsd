BZh91AY&SY��8� X_�Py���������P^�;"p�@ �O)�56S�iPj4��@ h 4�i�J  � 4 i�  j)6�&�hmM@   d�L�1�2`� 4a�h�!6��mS&�f� h)�<�ri�I"%D �����(��D�l%ē"D�r|��~r	5�408�w)�AU��a��k�ֹu)w���� �-,��;�7��9�r��i�h��!����4ۄʌ�q�s��`�F�NҔKf�\���ky�f�
�p�0B�`kW��J��x�[�����$�<������B/X�)_X2p�,X<8E��
��=��Q����M0��!�L:��)�x����(���;lq3��cz(Ѥӝ³�n�I��PX���2�qZ$�JҸ��p�
Zu�ł�@Z��(�0��Z	���X���&텝, \%����B���HQ�!�<�(��UX2J(�����\����.GEqYWVUe���.�Z�P�hr�;�c�1s)(0�%��
2ŖS6M�t�&��k��5���B)cޜ��pxLf���u�^�=e�%��Ix�������b4w�"Q���fEYବ���I���pdD��Ս1��g ��a�O`dC9�y�Y�Ġ{��Ai�y�Kg�2�^_8TG�K�5A��T*&o`m_풚bd3"��{�$���[]�Q��'^�1f�ɐ���85D�Apg:i:LF��Υ�W�7�ۃBrl0nM]���d���ϐ\�p���Qq���4�)��C��)�Z`Ľ	/I$s�7���8 �T�r	J�EC� H�2�1��IZ`�d(�CbJ��&f^YƵ�-�Pѝhi]w	{��:
����e@��t�X���04�	�������#BS 	��L�Ұ�D0?$Q"�xNl�`Ap�B��iTM��b��O*k�}���
��N�AHb<��`��17�B ��v��n%y��Ƅϣ��t�$�#���8�h�J�4�yb�,u�������£i�9��HcJ�$Lq�Y�G�2��@��� �p���MI߇1A*�	 �13��jn5/��Au�K�Ij�$J� $�j�c�S�H������h;�:x��ԤX�6`TRD�@w�\��7�Z�1�
��e���ܑN$(-N% 