BZh91AY&SYp.�� �߀Px����������`��w�Ps`
4 �J)�'ꟊ�F҃&�P�M4@@�@$��4�  d   ��⦏�H �d      Jb���O�@�� � 4� � �`�2��H�)��e0LD�3i��!��&Nb`�� � PI+����|�Z��&�I��M��SB�B�2�!&�-JJ!��>ͦ��8hD:+�i��`0IQBP(5e�$��#'�����p�Z��UFS]��Os�d��n��iSnpN8ݿz��x���i�1rEe[�$^��F����V)(�j��S�,�Pb��s�V��@%@�/�L�@3�+b��%_}��'%�Ĉ�����uQ�2�o+ ���*n[�wn�ܽ�V]���GG�_�N6�g	�rVh�arH�hu�e�X�MVЋ�+�"8E���T� �#E���	��
�U���m2���Zٕdہ�;�/]3Z��!$5|���e�YҖj��Ζ�6)�pEX9@��#CM*�<c�ih��b=�BҳK�8��<�!��-D����b����DXUm��:e��+�te���^��\ʦ{%�Vq�M�5�7QZ,�Z���NM�h>.�vj�:�Ic�h��֭ebҹ��8�����ᱍ�oCm���Dr���o��8��J	$:G+L�݌������d#"hH[ۗr��DX��HPD��Z�LLm�����+�Ub0�*�l��>
� �$I�[�/��双��g��9�f`������u��4a	:z�.�s�������RS�I���"�)j�c�� ʞ�5�j��M��A���o	>&�������r���^����4�?��'�~��*�d.�Q�K�"t���f��+�@GRH8#C5f���4��|�w��A�3w$���\�b��<�#����n�A�����|�5D�Q����L��)XR��tי|:�����6��i'�8i}��˵Fc1@L�ȧ�=?�r�J������2k�I.Gg]q�	j�M.iMR�Uc���c���HjL#�[�L��&k��k`��X�=��r�k�F�i X�� �>��x�������@i�\m��AA���`�Nf!Xnz&�$$+�GT@�Ņ�(64��ƨ�3]&755:��*,���"9����b�Nt�v���`H�z�l�楂 ���F��(X�����HЙn���$ 1Hh��ѭ$��&|�W:��0t�1�]�TmxT߼� �|K(�Pzc��׷~�%[�}�h7�E��&�D�T�C �A�9�0�M��`��b�X�Z�H�n��d3��#,Z�sH����5���Y#���a| ڑ2�lفPYIn��ՙ��mT��~�ȸ��
0�]��BA����