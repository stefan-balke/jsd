BZh91AY&SY��� Y_�Px���������P^�n݈qƍ 	D������H�44�OP�  F��J  �     BBT�S��yOI�z�� �P0`��`ѐ��&��D��M4������S�=OP �A驵<����@$�$�P //�r1K�LXj&�I����ٷ�d%�вd�&��UJF�@���;�����6[}u��3��[y$���`s��ϊ�b���ܴ���q���|��f̨ʗ;#�0N��L�Yb[.'�~��OC�`!V���*�n�IBI}aԊ��?��ƈ��
.�]X��AD�L�����	�<��\�qa��Oy$27�r?�h�WG1;�����
�����A���-y�'������Z�����YL��ĨU�h\=� �HЕQt!u� ����zU�\!��IlE�]D�q �"�EW �T�V�WZ��}�($�(�D`�246'��61���[m��m횸��In�G*���D�D���	&9E�j�7$lc�d�P��Q�g�$q2�-P3�eJ���k���	�6-�Xs2�ݔ�'��|���hx����"���L��Z��~ڈψ����۽���Kx]��@��f�W���B00`��ɿ�?�2!QH1H`u>Ӌ!L;A���pK_*���i/K�ޒ���5s�m<�EXFm"��jD����;�2<J�zl	R���KY�wx�&D\���-]&\�h��P�"�����aN�>�����K�C����Мk,Z6�B��� z���I�+ �.�>͙d�4�T�XIu�G%��N�^d�T9A�B�P��R�c��z4�!,%�~�o�ݜX�R\�ⶰ  #A��6���V�ᘷ�CFKT[k�%��� ��S�zv�����"�I0Ł9�����I1%�� Q��A(x�\���a.�p�+���`�#F�a,�nE�=Ky��B{k�%�r��̎�T�=gE�hxi3;@s�A��f�#�����2�Y�*H�!n]n��	�3�%qS��-�t���Pm9 g/ �e�!�J�@��7���v�RLu�udT�kq8��U0��!�V!�jzkq@䢺��j4��%t+� �����OW�'I��x:3&05�"��y@2� ���ݡ��f�m�j��v'��?�w$S�		Hq~ 