BZh91AY&SY�>�/ !߀Px���������`�y��0c�6�@V���Si����4�  �M�
J4 �      ���a2dɑ��4�# C ��MS�yM�D=OP=M  `LM&L�LM2100I"eO52b0��$��ځ������|��HZ�S�R�+���G%�0ШH��MT���$�4,�2� ;��JD%�O��q��x�w���1�����K7l�w%Q����c�Øo<��2�����l��i���2ΘۮUώ��/���*��ig٘x=-������k��c�������^��NK �3Gw๽�VI!o�kK�qisgP�@��f)W=�u��p����_CXfa2*l���9\�q�.����e�5��n�6����7PyXvfSq��ע��TU��/�_��:7T���ALj�$�y�qjwޯm�!��Һn*{6�6�*����t1SUh�P�*�Z����aj����2C��A5Aب(2�B�Ɯɒ��k���k)�CL�O�!4��)n/Q� �i��z@˧�ɧ!��T��L�2& AM�!���yA�f�l��2�����+�U�
�3�iˡ"����|Akx�j�Qf��'w]���� �k�(��7E�`ʧG{�� ��l=m��5�4�ؠ��=ᱍ�o�m���H�;�������#��@��͊��r�6�0Ī"#M��b�#�d��#UI=, ����A����RHb���H��a���P�iPP0�O���a	�d���K���vyZ�Jk��Tn���FR�ã���V� ���#f*��/n�#D�
p�=���"5����T�9�O�H� �{�٭��4ƻ)SF�%�A>��-�N�q�[�=pz;�?u�Bƣ'�^�lK������<��S�S�O.�`zT��$yF�t���d��3��^�P����{{�e�,tȟ�cێI�� x/=��P��r�:'SW e����M	3�E���|EXS��7!����'�v���m����3a �pY������YSZ�0��wy�ٲQI#��K:��_q�μ<�x/Zm�|lv����8�����c�)�%��²H�4i���]J׆z�3UH�noI]��Qɏb�UF��wYϩ��	0PԼ�PR���-U�����|I2�
<\�Ab��$$#@~�E�AXSr����/�T`x0	k�k�w99�����#�ė�j{5D\�y���=����Xr�,��{"jw\��b�S7[���t�+��J�:�8,uwnI�������;���d��8���R��8�R�*Fj�\��h#-���M�<9�F4������]Y�qfI4\��Y��9��-ˇU��ؠ�F�/\"���9Wҭ��j�ڝ5%�Y���g��1tM ��a��ъ����њ^H�&�[��(���"�(HIA��