BZh91AY&SY`B�& _߀Px���������P~�LC8di�Q���)����Pz�@h�� � 4ЍP@      ����54i�F�P��i��F�0&&�	�&L�&	�����bLɊ�M'�z�1� ѓ�if��RH�$�!�%��w����Q�
���P����]��Z ̰�h�j�#$f@���8�m䭧#��+�{g6t�i�N���Ó�ae�D��v�jv�4����c���>����(/���QX��"�l'���'%E6B	�o��" �h��HC���Ǝ"1�����q�1��eTAEUEغ�p�	�T�HK���g�U����]}��]A�Eƻ���tk�~��L,Dь‰��DP��W���u"B�TQ`2II��ق�.i9ZՒ���K��P��(�w��n��TX]19J�"�.��I*�)P (��$�{^�)i���ِ��ųH�*��&ᱍ�o���hi(C�����R]<�r�I;�ډR�/g���#�����F�n��z���G��Gh����Z�iAb�
�}���*����g��U��.��sk�v�,A�����\"XJ<�!KG��Ӳp��q�ԅo
k���25L7�h�w�tg�^�v��^Ѷ��.��3/$�}]:g������pϵI?�б�����=	fc������2n��2�$���2�R���M�	N7����#*Z�؞��BfD��p�c;�6'�����#�P�dE���nj�2�;i��Q���U�z��;2�e=�Fvɣ�dTJ�;^�#�z�¸�t�vv��`�1f�'��a��(��+��Vo-<��V1����3��̳v1Q��BZ�m�&K��Ðax)G���
�m� "_C�
,X���Ү|qǻ���6T��)=]ϘTx��U�7`hxͻ/�1P��k�k!�ݻ����@ Q��PE�;�X���A<0����eĖ0Y��Ɉ[5-b�xm>~1+v	;_!�S[�Y.�|o���kt��ǋ�gK�y�iM�뫴ܨ�Ǳ�u/$���*;
(���	10�3�l�d���bg�bj0UJ�
uu.�C
�]X��x[�%7t�֘��z�ӏ4d��M5�`K��$�e�j4�Y54�83�hӡs>uI�a}-2�Qr��K�T����RT=�;<m��C|�d�41oq�c��MT�fg�)�P-��y���"�(H0!\ 