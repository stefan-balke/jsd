BZh91AY&SYW��� �߀Px���������P��up�t4kM �B'�oT��~���  �@  �@�=@       $$EO�'�z�=4�I��z�  � s F	�0M`�L$H"d56�ƍS����'��h23)��%��Cؐ(B�b����YShG� ��R`E
k�s]��`!�b��G+T�H$c d��x3����xY�|[&�q���ܦQ9���Z޷���*f��uf���`P�W�@����g�VT@1"��r�=���m�uZ�]5��X�X�� K:�^�B�4,�����C��Y6��C+��+�("6�NOwHp��dX��m���yF-&�V��Т�J|�k)�XN�C2�fU�̰C@pj�D�d�]x9$���.�ҕ��`�D�1�2a�:��P����c(1�ՠhK3�N��V!��K�I���p�%D�4�1)"��ND$�C2 ��R��]����`�U0AQ�R�rr��Ct��x�m�Ӏlcc�m��Ar�=���[vʅ w��%J$%�0RF�#l:1)����ؽ6AԒ�(bi����,eJ���5�^�Lbm+������-��m��ߠ���oI]�`�oa~wgٜ��|�(�%���/)K�7w�xv��i���&m>Ǡ��b�m�,��H? �۳�w{��{��"ޱ�>a 3��c��/�)���РXP%�2
�_Q�lIq�B=�(��O��A3SJ�
h�bP<},��gޒy��l����Z�K۱�hdE�ٚij�qjLGIC�E���īd)أ�gGԳ2��E�
���4Y�]�� z�r�!i���(K����L0L��CNI.�H�7t׼-�Y25CB����N�I@�8�8�
_�T�Q�%�L�"/\q���k�W*2��$�WP����r����c@��g,%�
���39��XnxNQ�� �@9���|%�	�{�t��AX3|f#�*B!���*���Հ���<y47Dp
Dވ���`�Wcxd���0.��p�����m7���@��΁�h1�F�Bh&q�d,7e��]T�1�� f�E��^R,9�#s~pѽ��V[�e��l�E��Ry.�( �t� �4VP�jj((��i ����),�QXKڧ��L��z���&�� ��b04��a�\TFY"{ >�/mf�K-�3��`в3)����H�

�02 