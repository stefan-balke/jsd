BZh91AY&SY}P�� �_�Px���������`�<N��`{�� !��Q�'�A��4d4d@4D��0�h �� ���JzM�h4 4 ��	OQ&#I��i�=M�OP��4 ���a2dɑ��4�# C T�hA0�aML���M�� �y��5�+Et�-"I��4I"�W���+�$�2��J��
aS����Uc�t#CbL ��TJL�Dbd4�{Q����x�����&ݾY�r�2�ÌN��<A�J'��};k�x��HrK4���9r��Vm�K~��y곯�]�ڛ6U���Cz�[��`�+�cj�׺vM�{�o�u��$3Ӳ׺I23���Ƒ)A�U*`��*�""�N_V��@�Ea_pxs�5�b��Z�=u'dM
b	FC����DK��!�@P�[MS�K�����B��10���RrY;P�\��d% �6�N�M��$B18���	�"�f�;lZa�$E��&Z�R�h*���aW���V�ű���ET�[`�`oS���M��75Q"^�,&q����k�1E���0\�\b��s�ߖ,hpO�F�(�7˕�T¢X��G��H˗�(H"B�&�x�AB����vd\���ev�L�tI�Q��6�V�G)��f��l����g`�(��UX $���?t>*���%���i�(��&mci����D��"4I>��)'[�4�ʪT�F�bQbP�q,%�CU[4PP!,w] �H�>����3��3����GIs��b��ɠ!׹��+�m���@��3�V��R�6W�������D%2��T�݀�))�e�M\0~�"������o�?��?�������-Χ�}�[��)���ŘC}��}6!��jg�$����I8��No<�R�P�?\��"��'�|L��Jٛ"��}dʒ��d:�:��:�p���V�S)�(�"SЋ�5[�U����~2'��0tF��E�����LN�f^J��r���F���Xɡc�~?�[�J(���ؼ��������h��u�8�V���%�˳���.�.�)�鳻����ٿc�F����,X�T��տ,����J��m�\-̇����j�8bjx[�4�j�6ԅ��ej��ڼ�ְ�f��ȹ���+]k-e�C�[14�ʜ��W�vLc
����Bץ�[_-�Ow8��=n�&"�_f�#�u�����|746���.~�r�Sk�z��D�^���3a�@���(���Cqt.��Y�O���֍>�1UJ�)���b��Z0U����2S��I��-GMRM����|��+N��$2j�e����:�j��'6GL�ui`hФ<�n�L�F7��K�ԍ�J�ʤ�=�;<4;���je!���K�����s���9&�A�'�ߝ��w$S�	� 