BZh91AY&SY�2�� �_�Px���������P�q��8
d HH�O�=	�='�mCѨz���x�Ɉѵ����)F       )��oMPh�<�@�  M 9�#� �&���0F&$	1�S��#����OI�0&����� �!"�����P8AV�$�S&���m��0A�hW�]�A�Q2��V�Ʈ�Z�.�T{�G�Cߥద��6�H�x�u��j�b����:�"ISQ�Yb�[`��+?ފ��d�[�+�.1��`�k'1�VWJȎUc��E��!�\�;��BV�|ɂB�Bz�(�1�Nu?��V.��$0�Ɇ���c�ȹg!]�AtX��ɘ�^>�(.�+k�䘛b�O$�>�C$�����]"�@��k�B8�PHC����¹	 � �O($69�b�y�Y�{("�*��eG���QIC���x8W�9��������]X����$��h����J��-��W��UK(���t��Eo@E�TL8��I`����e����!	K�$�P(���`����p�4�������+[���&��KbCm$P�A5�&�h��������F(KfR�! �����3fC2\�q{xnv���G%�i�5m
��guw�8�.%<�e����/"q��t�~z�`Qc�%����}�{�I��pkfe��7x|R]����|�	��
�-��v��B��0�_�2��/?Z1�c�<ѩ�:ͬ��4�2�@�{"�i'��*��i�����tj��5L�P�=��� �.��C9�L���aJ��ă��C��4,gY�mƒ����^��������Ҽ�
AR}�p~_�5jL��q�l	��H�:}U���8�	l�*�!^ޛ�J�P��2pb_�~K�r9,�\$g�:ɠ���W�A��V��ݵֆ��H��=�4}zG��k�^s���oJ�A0�P��Y�MT��H 4�I�8d
�+]�llj�:��b$��ʓD4T=�@Q6D`mҏn�'���GI���vt)G����͆!�����#i�{Q�j7�>��hL���X�H|�h��1�{6�B�L?�+1c��."��T1
�4��$@1Q�$8�6��5�߈����g7�E��&��f��Q"�� � �1X�P,p!m7.�a��6a��),qR���
�ޥ��4z=��&#�A�9�d+� �q�فT��7����sk�ީk�,�4lO]���ܑN$)��� 