BZh91AY&SY� ! (߀Px���������P��2�Xm� �J"��?F��xSC�P=�@hѦ� sbh0�2d��`�i���!�HD"Hzi=M�2�  �m 0&&�	�&L�&	����LɠM4A��  z'��KI'֐�BH�h^��T ~��ts!/� �B�0E�L��Ŷ�xX�hZC4� ��5N�ARﻰ�������wZoNɔv���xM+ڣFi��$�mX�C�B�.m��D�	�^����{z�-�H�ʍ��]i�֘\3��)�N^��N�d� We�Nh�+F�oD�0��an��_)J|<���Ð��;s�����иn/w��m�1�<�Y�e(!V�-7EL5ቺz�����oG�X�[�K.�` ����PZiX�rr�M�QYY�����0��G��V30�3l�j�ф�m��v�Id���b۪�;œD�����8�	�!�=1d�T� �d|Z-��Y�Y�q�\vf��,���5�9+���k؅N^m��)n�V5�r�Ȼ%��r˱��h���>���A���o���hi
���gp|T�i�R��(�(��,N�Rt5�(�k7$lf�������6䆚G���@ހ��AA@�5�q|�Hb���*jd�U��fIc�%���c�����_M��`�ܔ�\��)�X�S�/'	�a�4I"�V븕|Zm�7)���g�sb��Qot�"B��>rʫL9p
���B#�A4	�yD�
A� ���佭BǊ�Vԗ����%�^��4������h��+��� �I��{ @��w���ҕW5�emYը������!���2inipMg��3d'˂��=��e��PC>ºH�ʂP��z �-�|f�Sp�)H�`H7���=z�!t�i�+2(�Du�A^[�D��8�&���e�E�`�|	A��aј]�W�I�1��lJ ���`\=t�;��CJ��@��7_Wy����h��fA�Eu����,9������E��-8�^�PY��$$#�I$`7�:�ْ�2�J[$	ǫ�ͨO���H^|��"G�|*�l.�ǲFh���؏�5	��9���)	���i��@`Ύ��-A4)g��iY�L�9
�t�cM9 g"1�M�,H�l7��{� �X��F��э�{��LY7���� �5u�
����s'ঁ��D4��G�H��灱��^$]&!���J�����6�|wZ��T��f���`д\wW?�]��BB�T �