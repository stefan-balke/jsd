BZh91AY&SYl��� �߀Px���������P�e�g�F�!(�=S��S�=���@� �jz#CR��#@      HH"e
4yOM�oT��=OP�Ȁ9�#� �&���0F&
�@�&i�M�jz�H�=L@� �M� O�BHAt�e$���z���i#��0Щ4���b�ٷF��̰�4y���H́���u���+�Ο���\ �l[�(��?����j�5n��U
�-~¢W�T��o!��9��^��L(�L��C��=�ǰdU�d�n��v�`|��B�[��k�%�MU��۞��{69ˡ�QUQE�]xC&6!2Ba/�R�JW-*�}�S��^��0F�1���r"h͜��sPn������B4p �3����� ��Rk�<�B�K�ȭJ���Vhe�$�.Q� �� ��	T�$��͙Ig�X D�!pRP$�%���7F3J��PED��J*�)	�jşj����ʳ�=fj�K�����m��y��g�%%��#�
�>*%J$���HF�F�H�(�aX K���ӶU6AIVXda����J���k�%��1��pk�rS�~�ݦ;G�Uo���O�^b7�0a[��O]���?5�ϗ�RՀ��t��Q�������F1��ש�=�5�[5��#�:z������[�xH��Q�hX�hwW�n��y�R��M�ɯ�N:Q��?�2�$�h�#ȏtk����
���K�����xR�?�]�JӁv8�RS5#k�cC*�n��ܳۍLLuʝT��{ec1[*w3��e�Ȕ3�����%�PU��M[̌{������63;&)y����~�f�(�<��N��ٌj��f�ҽi�����n�F���/zW��CE8,
6��4��P�TA��d�� ��h�:�Q�4��ǁ���Tv2�WuQ�;�k��wL1PԼ�R/����W��j_(
;=�PX��%�	�>�^F1v4�J��ح���b�k�Ert�����[���$�S[�\����=���|�ѱ��Xr򳋮|�mky^��ި�ǵ��2]\��Tv������{������f7����U+<)�Թb��]��3�Gqd��y�+FZ:$�q��K`,��ì�#
#pg�n�����.lˌ�R<�.�f�Uz��"��}p��(���nM�z�s&靌�{��6;��mz��|��3�h<C��7>/���"�(H6[B� 