BZh91AY&SY��� _�Px���������P��]i��dր����
lD���4  �h�L�����   @!"&����=&MP4� !�9�#� �&���0F&
� ��24h�M�򟨚dѡ� Pdф�W\�-F0L�B���WrILA�B�`�P!M~�~ 8��`�бb� h��:	,d���s�v���]%�����*�b�W�,?3�-�nWX�
��n�6�
�m� ���Ή
�'���_q-�!"���g5��BN��%C'AK�F6�77�#qjz{ ͵���@�!L7у��2+:I���L��<_i�l\:bi��n���g�]j䥧SՃ�U�Sk�%�2�Y�`�<�8#*m��xF�r��E2S��L.�͡eJS�H�P1h���9C���j�/~8�P)����+i ��Z�aa6�ꮕ5�^ŪM#S�`�lTi�O(s&�#��ӄ�0��]�Yr���j�Y���Z�,�ӊ��!�h˙�>f�"���a��}�6��\[z���f�2R�D0�/�61���m��B�6q���᤹8H�B���~�R�-V/S��j������cM�(�j�m�aMYPA�M#��e�[*

��Ku��3)�M�0��x2�>1�)��Ppx�y{XT��%�DMv_��h�y�����!=XO��؊�w��jŶC�۔Ƹs4u�A�M
����wp�=��{N	5s��-���9��LAKC+��{􉷶�g�$�y���pD�F�t?�LR��tO��R�����̄9�v$���a�9̷1M�����m��ih�~�-�S����S�.��X'+8Hpg��в����K���f_�cY[��f���u�='���f�E"v�RśV���������j���clhd���U��v����q����6��שA`�$�� &Zk	F�8��z�2'T2P��r'���*;Y|*�6�q���l�ꑒ��-$�1���ن�/��"�B�ƽ�PX��Ą�b^�Qt��q�ܦj�L"�#"KaJ+w4>>�&��bف�b�'H���vW�m%E��÷�f�Y膷���9���;݆kȕ�X��(�y�"l0��ݲq3x�G�;�9LR��;;X�]��*�����)ѻ"e�x�C~��ߪ��da/\zv1D��u�e�9'!�����߉����TN�7�Q�.l��_�R66{�v�MIROb��+�����3��Nkŝ]v<w�̳��+��b��V02������)�h��