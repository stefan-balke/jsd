BZh91AY&SY�`  )_�Px���������`�<sa��t�����4=F�Q���@2  4 J��T 4      `�1 �&	�!��L��������2��&z�Tт�z 2�9�#� �&���0F&
�M	11O"����MOS4�1��e5/+�!i c$�9	d+����ZH�2��EH�L*)�ު���!dhXC0�$�<mU"4H�1 e��|xx_��^u���ܜ�=���z3���'����8�:,��~��U��{�T�3(�qK���3�4<(ho�h�~���9�
s'Q�m���F��*JT�!��;;_����tk�kU^�B+N�\����F	D4k�9���n��ſ��3�:t�K� �=�_ ����v��۝+�StE>9*/m���V�rО�e�xL��H61�(.\�\�Kf�|L�-KZo�A%���e�VC@n��X�O��m�b��:|#2���Ec�Q|G((�RV�[M�Q���L".8&e�q���Ա��3,Qj��
,����W"�����5%�R3JH���ef �,�`���d�V*�.B-ziN�q���#<�J�w'mY�P��0��{�,K�mT�N��I|�U��j�ƌ�y�g/T2VBT���s&��TI5�ۢ���C�w��:�bia�|������m!'�w�A��\���B���D�D���k�i�QD�V��#j�F6��(c��1��FS˴�4j��IB٠��a�n����u7����]9���.���*3�ꖢ<(2�Ixj��.��P��%pY5��mtO#]��{�7)+K̍�%����\�9�I&�9�'W�	x��}�w/D�����=17(G�Z6��+�߫z\���:����F�	�|����L��T"�{�m8<q1JvP�=�ļZ�؟W��Y�3�{�4c߂Z4�6���|�����F,<4۝LH�(���$S�Eʚ|�2�����S�-qVS��ͲutK"�U�1;��e{¹i�n�Zf)c&��?\wn�P��'��;r��.^�GK�o�*1��7ן3��.�Wr)�������ѿw[���=s�DX�ms��ԭ�e���"��l���>B>��@��e�W�To���6�fÜ(l\먋ݸ��W�|-�y"j,,QǡA 櫓!!�$.�p�5�2V2엋Tdz�"-zZŵvm�zyD���-�>Wt�M�V�L
G��3���k,;�vqr��I���W�y�y^gq�E|CaR�k��F��]��:��ϕ��M�U*U�N��0R�cV�m(j�6Jo��Zeh�I�L��w<�7��뀐,Q�a���p�Vk)��GV�y��8m6&(Q��F�=��#g»68Ԕ��Y��o:���.��53�݄Y϶Ƿ�UT�9�s���r��ED�0u���"�(HQ�  