BZh91AY&SY�2� ߀Px���������P�;���h���l���SiF� h�  IO!I��Ѡ�H     !!
dMC�a4  � 0&&�	�&L�&	����L@��ɢ&�$��1 h��zO)~Ni'�!�� �?�u�
&,5�+e5�>�m�}��hY3&4w�R1R���n������^]���*ަQ>�N{�ǳG�D\��P�-�~�<G� ym�9Yi��8����#�Z�z�ۍz��#R��� I��R@*���d>bDC�=�I��L:D4���?�H{����w�B�ȹ쁁�{ʙ)�G��t������4����0��XȇM��72�jh�FO6f��2�2�cy`z^�$����/��F��aw�ȃ5��Ǫ�5#2�o<�\1���;��HC6sq���o6�m��B���⤹��B��9h�(������ڒ7$le�?�FL�F��ƚG ʨQiE�
ռ�0"k�9 �<煔c�d�s��@�8�:yvS�����T�n�=2����<p`� �چ�D����U����8��|C�>A�+9�!���/:�q����z��������F|��2��/I�vD0���l��	�4Ak[�ԗ���32a��dx��I<Y0�����Vљլ���6�2�������D�����T8���A�n(p3���^lX]9t
�����dhjB�&>Ѽ^r�}00�.Z㢦���N`�-Ĉ2�'T��v����+X���F�e�y6�Գ-x���q/<���I]}��!���	#:oo��R�#��L.9�Ve[A��k
Cr�*�H����PX��%�	��%�&�Tf�+�P�!���PI���nByO`������0P�zU0����@��34��u�6	��:�YRC�Ѹ9B��k	"d�=j�³�� /���ci�8��T1�p��
�#y1���
v"ujc���0��\�B&U�8��ƠW&�(�[u�A]cG):��41~�.�����kI�� ��6��QY����T�4���h�]���5CB�����rE8P��2�