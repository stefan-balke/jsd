BZh91AY&SY���t '_�Px����������P��� ��2��]����G�jmCLCA�  � %4&���4      !"j�z�'�� d�  h�L�1�2`� 4a��b&��=��2'��'��S@ bi���pW1$�%�LB����Y��/�A�B�0E�)����n�d�4,!�a h�j��A����n޿,

5h��T�jk�5j��q6]8��+4��t����+�����F����w��J�
���)�.""�9!=J��2�K=�9
�Y^��0Zk����r����y$a��_A�q��6�cw	p˗���U\6&a��d+ud�q �N�#n������$T#-���S@Dwɔ�fi�ieؾ�D��X�6�8�ۻ� a1�M�T̊�I��&���1R�I�YI�8��\�Xm���|����߅M�aU�3AzZИ��t&���ʛ�.QI�h���s)���1e{�-��c��ѥ�F�,C��=���� {2�݌Ғql˴��1��]>0+�;�����-�im�խ6{p����v9�cަ�m��P�v�C�:T.N"9P�'yݢT�K]��mT�2�m�/VD�ٌ���K$YƆ;AԒԅ�e��P4P�(((F�����Hm-<ڊ���O�\��3���1��ǧ=�^�}�Í�ymв��ݶ���3�
�|����B�8��Zm	҃��Ǥ�\�1�f�:��'�������N�a��$��T�����f�]v��ڗ�-l�j��.��S.N�z���;�O�k�O��ѝK9hm��g�Sk���K,��uI+]�k�Ѧ���ki�o�y�a�o�"\�i��]	��4-�%
�`֙|��F���������qu���(��#�yϸ�aԯ�l*�l
�ˌ��8�w�|�`L�a��!��f�&���˃2�WEF���n��-��M湞}l�!L~[7��8�b�D�ӌʒX����}��ߺ(q�wXG��D��zEG:�:��5��^c����.P�.1����b7m�=#@@ Q��A ��Ľ��E�@VL�b���4��a[=-bھ-���^����dO;�3�kq�eH�v��>�m���}no�H�nn���mTJa�z�3bJ�"Tq�ϺD�g���i`�zt��Ӊy�6@h8��DX{Ԍ�%���p��VC�@oW���KBι����P8�Y��R��6-Fi��͠�ե��D�n��J7l�����g�U�i���΃I��dp�di�n���t�^�^h��V;�j����vh�)�Pڢ�qb����"�(HI�u: 