BZh91AY&SYyA�n ߀Px���������P��@�d���F��D� ��h4  	"4FE0��Ҙ��4d   !"jh�F�C�hi�Mhh 0&&�	�&L�&	�����$���ړ�h�Q�bd�� h�M<���J�"-0��{�Ir��?%\؏�A�B����S]��|�f4,&a�8�D�������j�u,��蛦�r�D���n��o%���E��n��mؽWR]��$o5~Y�H�kH��P��h��a˦�l��N�͙�S�#%���LEq���o�F�㟩ш+�����q�lv�9C��ъ�[_�K^q�e���:~u�Jm�q��6.�k��<̌��Z"�d�*�	�5D�80�$�X�)�3gq��WQ�Zei*�xL\�F��2�N�L�-M�h�*�ʙE�w
��y�"���t�e��z�N�8��������m"��5���#�
C��T�Ix�\���]���ԑ��":&P���H�2�^�gD-�#]�S�0�kSO�U7�圚1�h�֝��Q���a7���f^'�],�?���
j�fek??�l�cW	ŷ�SI�h��2ոQb�9N�i�����5u)�б���^��|�y�R��p��~����p�wwvH���Κ>X%<44��_��0>��Yg��2I���)��6��ƻ�`�ͬ: �Z�(C.���8�LY⎥A���Χ��ɲrv,�l�:421�+�6�ÓCsS9zX�wc�~��(�y.7��:��c=8�M[�/Y�дc~4��2a9͒��{�S�߳����5oݱ�:<&��,[�whkV��=�<1Q�m�#\Q��y�G��̮��Lmf{Y.�b��y���یmU~w�m��-D:���|��	��%�.����3@�b���d
Y����s��%i���`)�Ӛ.z�G}��G�73Sap��l���Y��eu�ʉL:�;��t���G��=�f_�����n���5ubr�*�_
tx��JL*�r�ȿ�Pcn�2�ic3Jȩ:ԛo EHq�sa��f�	@�m� �UO��s.s]Leݕ#o}n��*L��Ο*󒆑s&���6�78q���媟��Eq����hIၐ����ܑN$Pp�