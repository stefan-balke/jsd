BZh91AY&SY��D .߀Px���������Ps�3b�4 Sj&h�zOSj �     %L���MS@�@     		M5�i�4ɰ�h�   ��b�LFCC �#	2�50Ҟ��C� ���)���BD$
�d����G#@�8AV�!��&I��_)����B�hVf4s5N��3��M�86o�z�޽�+g�*e���`��b���a��[E�mڴ�%�Q>��2���8�/ז�����Ac'0Â03j������ V�<ɠB��Cc3)�|e�Ġo�<ڼ7�t"��p��ZYl�s都��K�ڻ��|3B4/�LG+�&�$fix��:�8��6F����	A�b�E����L-��'$aZKs,5
CEQ-�6��A�Q�Ac�H�0�Tiȅf���y�L��z:.���C�g�Tam� ���7�m��Сn����%�a�R�n�R�%��dX����#c>�r,[��x��vXd0��	�"A asgfLcHm���Lo�
#�|ĽaB�@4�#.�o�!� �eA1��Z�ǃ� �����a�	���n錣�V�x	�m0�d!}�ٗJ���^�*o/�B9�����,A$f��Ќ���2�)/N�Q����:���bc@�fE��� �-Ғzh�m���h�:�in�C��+VS��!�:���"`��Me��b;��mp3˘����4��\`�i�Gx��~��\j] �>��?�����K��8�Nj��n��2�))�d��m(��3�����O���f�V���LP�zd�־ݻhд�Z��^�i�G^q�6P/9C�EF�K�j
�s�r�	�,�#�R�v�`HHF/I,�`��8�\x`&�h�w��`��>�'��א.s�Pbwb"C�.�݉�� ���F�q�X�@k)��8�Đ� PѼÕu��M=1W9Γ0�E�@�N���!�Tp�/}���̶n�*�+xn�i7ZE���ԝ��
�|�A�g4&ơҁ��k�Xh�)-0@�F2�)u��=^��&����y�\��D�
򢩌�#�t�u�^G
���h24+�y����"�(HCl" 