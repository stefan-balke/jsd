BZh91AY&SY��F� �_�Px����������P��9p�&�0�Jb`j��P� � h 4�5S�h�� d       ��4�FS&����P=OP $ s F	�0M`�L$��LJy5=G����H4 L�W�WT�I0�H�B�~��W9��D4*���5����{,$�4,�����tHā�����;���}ZAu;��/^jf�����]/��|�H��v�C�.��� %/k1�'����0�A���� nMp��pVd�$��G��A�s>Wk	!c�Su�K�5��D����d�k��[�|z.��1���}�����]��˞s�]J�M�y�S����+$�qZ����f��\e��T��Q�
1���h]j���Kji��rkqa�1�MKT�n��4e��XfU�-�*eci������s/W�	���ntꭝ�Ԙŋ44��$�� �KXᬘЕ�� P�Ah0֞��_[iKw&���\�z׫�����[m����;lq���wzH�B���D�D�t��Lh����b�֒7$m`�i����2F�[PP0�mؼ��&e#/�My�GC�G!��uF<�H�lGO���6�8�:���ˀ3��J}K@>`�}c�4*��%�Q�j�Z�gU�8��o�_$
 �!�N���/I�[�yI��A�����K��6�ڗ�b�����|4����t�=���J��M�v��j��.�ۦ)jm`z<)e��\����q�79�Ef��,�Y���j�5t�]#��S@2��`���Iv+xೲ�b�����T��dRJ�]��׸�eޯ�����3�L���������K��eY�i�tu�'ǎ�6�%�7b�D7�HP�lu�+A����&�~ū�g$��@%�X��N�V�LQE�R�2S�I6c�<���ǽ]Uu����ve�21P�^j�_{���W��j_$�V.q�("����$$#�]"ᐭ�S%_{�j�O;-}(������l�T/��j����9^��1a��s��V����t*%0�|n&K���j�Q�R�:����	����������N�b�T��WR�)C
�\�h&���M���&6�ttCS�W2_�|����`�])cc�sU-82ϙq�J����Va
5�5��wԎ�p�o�*'�g����Ct��7MI��޹��Ǫ�5S��e����@�`d)'.��w$S�	
Th`