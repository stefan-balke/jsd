BZh91AY&SY���[ �_�Px���������P���FT1�&��V��(�2i3�!�i�ѐh�h �&���P       HH$�$��OSQ�ѐ ��40&&�	�&L�&	�����(ɴL������zO)�OQ���<���%p�%��"FP,�|?��W9��� �B��,$2���f�;�6)�a h�5TFH́���u����k�+��6�Vg��/������r|��h��t�tç�pvi�C�~>������d�x���E�c(d�wD2$Q�dB��Z���Ky��!d4A�	��_�6M���z�h\�,!�L�
[�1l�b�W4�T��لI/g�)�֫2啨���%�.�Mj�o��E��Ga����zڎ�2&j�A�n: ]Ej#�u��,�ٳ
�n�"�d
AH��!�qHKj��+)2���̉�����Lu����*I�BKZ:J����ܻ����306�,D���2�^G`X-$�
M�nԢ�c5��d���0L��3Y7K�.ف�~�����7��m�4�|=�g�=4���G*��>*%J$��aq���/`���ܑ�62^���O�H]̰ʨ([J((96�ȡ �	3$4ڕ���vh��#f��3����ǏV�[���			�}7�^��5F`�@M���{�A��S.N.>E%2�A�=19�	��
�e�/ZH�|��N�������RG�Z34�k���Η�����<�����e�I��1�<<c]7?��47O�(�ũ���稜||�JՁv8�ɘ��R9�n[�P�2#��n{g��ˡv&.�B,m��U�}���83Ù��l�J��F�#�x��˸��ml�%�+�Oi�{�ٲQIW�OJ�Ռu���96�^�m���5%j�vy�y�/��jdh�;rG�F���bŹ���J�`Ʊ�o銍S:�m�zG��򊎦=j��p48��d��1P�y��K�l1�V�ٯ�iXXQ˂�(,A�Ą�`��V0�e���k`h��K2@�6�7��|Jۇ:Gc�/�ߘ\���+�=����;2ë�g�w���n
�:�qu�K����Qĥ�zR6Ƚ�l2wf������i�8�CWr.U�H��n���Ù1�c��s8es%��˫�G��F-K,�;[T�s*Z,Nk���F���b�GK(R����_H�ʶf�*I�,�����7H��t�ę�+���~d�Q[B�|ѬV9��a���j��H�
^۫`