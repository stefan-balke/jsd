BZh91AY&SY�2�� 5߀Px���������P8x@0ƍ4 ��OT�����M�=F���h2���&L�20�&�db``F�*z� mi���� 0&&�	�&L�&	�����O<�I����)���@�='���@>�"@�H��� |��ѭ#�bШhV�k�?6m�氅�Ю2�"h�*����2}�鳫��ٵ��v�n���pʙD���p�&+'5	�eJ���t��>T��Ž����i6�bf�b�$'�|� فZOQ�jӰF+��� V��9�B��"B�ȏ)J�����(A4�����A��Ҳ�,�.��[आ�'�s^/�5Iws�J��pnb[MQ��<�GHz&kfR-ToR��]Ѕqҡ؆����0�Ya�lm��� �da��f�D�g�X�x�<��`L�&�z 7�W�=/10�Wʖ.�x��z��T5Hњ4Fk�����m��!��l�%ǼG*'���*Q&�ۤ\����Hܜ��\��9�)��H�2���([*((F���hET%]M3�u�lo����0��N)��D�d�q�'�d��S�hn��4��K
W�j�8���U�{p�#����r��e�i��3�gdG��	���@�Z�!+@� L�4��.+�e�$���V h>�^h��ϕ"��kK���̠{�%�RO
�[T�]Iɋ#��c�Pf�E	r�85A2�l\!�,dgX�*�98n�Z�ѾCig�C�
Fa`�P� ��;Y��֨,	��Ju����+�I��A���F5GG*����� ��vCEiT,�Qٞ�hs)��C�)gd�g��3�/K2[TF����$�voچ�-ʻ�t��H�����P.=A�ķ��a�I���+�T��HZD
7:����2Ą�i{��F�%Vm5�h(X�!���*%d@E�u�n�'�2�8)���$19w�=�K� ���Oj��3@s�	��z�bHO�(h�aN�Z�b��i,z�Y�8�G*��A�恜8��lEbH��0����g�~"�"׆<��}�X�%:�)�7p(
���2z�/�\���o���$������J�j}�}-#�ۉ���xzy�bd�����H�v��6�&�Kh�2Ƣd0hR���O�]��BC,�^�