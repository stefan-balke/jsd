BZh91AY&SY�v[� }_�Py���������`�vˀ��ʂ��@��i�L��ɂ2 @ j��`�J �  @  2d�L&F@��M#4i��DI����    4���4�	��0#F�` A" ��P�)��&e� �"zMeB|B"�]	(>���rl�� �B��� L���F�u �\e�BI���rD	+�/���ᷜ�&�h�C��#�ܜ��&E&K�L�t���
��>-����p�3[��-B�2$�ڒ��ky��W��,��{j��E1��c��w�|�ٳU�&����-���*Us�%Ör[kË�F���<hH�(������KAe��f�:ֵ���~����'q`� "���-����3���b1.A��V�C~(�;�*Nb�N?
�����,. w��$&�H����Ƞ���/��Zێ�bEa�j�`�/(2�f�1]�#$b�!��D�n(#1}ljF��Yb�g� �{VD8RA1��Z�ԘL�'ۖ��'��lJ&a�f���xڵ�ظ�)]i����)�7,v¬F�*�F�cj��fq���k���d70�C#�	;��,��F�xg|i�)��|[F��a��S�Y��%A3M��X�D��X�Ʌ'@jgG&\Hx�Y)ʙ�fǄ�e��c_^�,
�u�t�B��t�%&�ġ֚�d�!Uz���uX�L���M�����Z����61����CHv���C町�Hq0L ��R9r7TU�a&�hY�+CjD%���i1��+1�����k!�D��I
��"�R`1���d$CYy��LhHm>�����ٝ����Nb�^;%�H�@c���n�ᣲ����	d�{w@�)5��e'z��9�6fBfa�y ����nC�EH��S�0j�k"��`1`в�yF����(3�?��؀��^�ޒ��IXB=B�&s
�D��U�t�&2�P��VAq~ē�P�Z�mE���@q�|���(4d"�te�Y ʡ;\I��5�+�^U/�t_Z��6�{@�
��.�	t�(-����(��f���y�@�$4%u���G-���M���T k�J�*!J�Dq�qp��K��A�M!� X�Z1j^:C�ַ����ƒK������4yu��iP��{K��q��؈
�p]�[�/iP h�bI���V������;D�n��uE��j�p�A)�٤�;w!=?��Y�%P��f$I�@��gxr�&&$�3{#�eÍ&�xB�PL�I�p��,H�b������ W
 (x�.u�!�t�aQ�聜8��J�"QA���A�to.3��~�ZmA�$�f��r�
)x����XfR2Hg�kCP�qP�\1���ƀ�+; ����E�ا��m��m�+I���1�b��@Is��Ȱ�L�7s�wsݵ�nU��3gf��ܑN$1ݖ��