BZh91AY&SY �$� �_�Px���������P�l�݃8�@�%5��O�F�5G�2SOSF�jzMSA�i���Ha�L4dh2 `��
4�� z54 # ��9�14L�2da0M4����$H��@��)�4�Q� ���zM���(I�I?���ZFÚH3E�(`$���|��9l�F�a��$��)H�@b�8���3��GO��t�n�����>��)=I��ﲜ�@��z:�3-��V���ޔ��Pؓ{�=}��8_	bF�����.�1x��zIB�����2Y�\�I,0n�B�!������6ʊ����_��|`��!a�y���s��&��ql8�BX���t":�LB~R�����0
g������kZMg$�[q��<�v�&`�Y�ňm��J�`Z��|�C�G����Ҵ���!�\��"K�ZdVUI�\ڤ`2��`��-T#Pa�t��\\Y{�}jke�)��pB(����ZY*�K=ʩ�0R\X�G�ʇjV(]��h����a�0ý�|�c!�-��Y���`s����lEwU���$��6w���pVQv0ҫ;*�̊i�42hjNZ�7V$j��$�bDQ�"�5D�W21��ICV"$�TPP ��P��$�0�G5#��z��r��W'Go=��� HG�s{�����<����Ɯ���U姄�
��Ր��]u�u�C=ɇ���b5_/F<�������x�����/�3�p�_�Ba�����n����1k�z�iA^A�3�Ý%�P�z�f����v���8�Z=.���T<~�� �-�6%JV�*�n;�naA����ǞAD����� �0j�JH�V/�!���%U���@�m�8�Ƨ9�0E�	�@������u���XS�I��>_u3��Do!w�GEQ��_�0��L��CE'D-�ٶ�v��ZcX��%�U�G��fJL�4d�!��6����Mv����ˀB5,씉{c�Oq� ��w�<��ac"�"Y��H��d�Nk0vm�T��I$
̴FjH(@�a1Ȉ!��H�E �Y�e�9��(�4X>b�c:����Y���)��v:�jy;m�fx�4yUl�����1��a�E�Ʌ�,��z�cHP��⅙�1j��k	��C�֮a�?��"��\&6��3�"D&N$��A�Е����`3~�2��n�GH�:�Ԟ7�PQ�C�p�����@��R����P�Z�A�RY�(�����ZF�����id}���F�&l\nE�j�n������I��B�tc��q`�5�-���b�H�
 d�@