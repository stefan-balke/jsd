BZh91AY&SYɓ�K _�Px����������P�7w[��p� I$�H�4)��S��'�&�@4���&LR@ h�    � JdBjj�4d4�4h4�  4 � �`�2��H�Ah4�JyP�т  �dу� y�B����?/o�9�aZ��M$� �^���n�4$\4+,a	���9(�E�s���嫟,�ّf�H���92�35�v�
�!�3�@�|�2���6�)BJY��<M�󭤐~�;Qn�Z#'���Z3�uQT��٠V9N�a\�y� �kz]� ��L�����F�S,�2}S�Ɏn���d��S��:2i��VHܮ=�H��]L�˩�%%���I1'.=�ބ�*Z��L :�< =z.�
�4��AȂ�P��b�J���hd��ZTR��&�Ap����S�nL	],2�slկ���%Q�
����P�a�2�p`D#Fe ��,U)$@�b�e�`�o9V��t�k4)4١"�;�hY%6Ɠk[B�YԬkd
i�R ��݁�FFDX�"鼂�D��#��	7z���5b�f���W��7��$!-��I@�3����I|#NY1
ϊG.F��IBI$$��t�4pә�rF%m+,��L���ÚJ��";H�E�3��! ��ߍz"��#^U����M/�f�T�q��Z1�����vdÈ�_�#T�Z����5��įo�3�N\l�P�gz/$l8Z��.  vcY��k_��?�l@)�$� pX2j�����r�y�'ߥyn���В_�53q�!��1A��%풢!�I�
��ŐA�]�$�P%Z�~%Sv����A�����|�j�2���0%���╅*��/ZP�3�дԯ�@�����T�Zu�`�]��K�����/�ޚ�@4���(k)���<�#�uw�"�CF�s(���aU��פ��19`�nYQzIo�^�8��W��������pVA�H~�]9`2=$5�r��@��0,#�(00&X��V��\�H�6o�HP�lP�lhP�X2ttL1*���"T� sd@F�~+��'��K�����
����lf��0D��9}7����ُ�m+���!a �RM�3��zIbJgy�֯-;��1ZwT.�N��1���q�B&<��3(3v��a�3�j3�E��Rw_ĢIT�DDM!�j&��[u����F�,0��P@bQF<��f�����ɤ�k=D����$�Xe6^TRD2���Z��;,��ј�уB�Io�.�p�!�'H�