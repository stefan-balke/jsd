BZh91AY&SY��� L_�Px���������P>�]Fô�j�@Q�?TzOI�$�Q��i��d 4�h�Dj�       ���)�hi��S�d��@@`�1 �&	�!��L���L&S�L����S@��5����@����Y���~c��/Af� Ĩ$�k�E}T��˘Bh�j\��E����ӆ�t�h+����L������jz��W���htr�9[&t��e������2�,\b9�`Azs1��2�K����-.s��먐+��G�B�w��r�N~���I�y7���v�E��c��#�/
����fX�3�d��b�!B��ilg�)HF\I��c�d,��H7E$��MK��P�.Y�(�3Z
a-��������Ud(�%!������[�ሡKإU�*]�T"�(�RI0:��6򼴌o�(j�X�LbᅶKf$w�c�v�m������5q��Rۉ&	I�<rDđ��sO��bŭI�E���%`�!���q6JF�Hɘ�AK�HH0���[�LhY�������[i��x��<�8x���M}#H>s[+���������1)7��~�[^wz��f�Ds��}�+Y�]&L��$���d���� h`��j�!A��qQP�@��0�����0ԊKOp)	y#6o<h5`o^VBd3q@��Y�i'�U��6mV�.C�f���E	�4p5T�Tp4p��f���m
l���
��(���.6��	6�N4(��
���������AR}���}-�`ĺ$&X	�qȿy����8�!�X�t(2�-� �L�&s/����1�.ݦF�/E�-��Zk
l9ΔvP�k�X���sH�tu����ΐ�ib\QQ���d������崢�@:4P"A2J�Ȃ ���H�^�5a�eI�* 6Dc����B{�K�s)�̏^@�1r�{{�#3��?��N!�Y���7	���p�Ĥ�h��N薐�S<�[���:EwUCRfAQ�ꁜ�!�*�D��c�Q��q�UȒ-�q�m8�"��Rw��PJ��L�`b�����\H-a��RYB��YˡK��fg�����h=�'I�/`pJE�
�i$A���̓h�8�Jݳ�f�A�`Я�����)�e޷�