BZh91AY&SY�� �_�Px����������P��۷ �Y4n��t$�	�4����4���@� 4�J�)�dh�  4    $""h�S�d~��H=M� h�h2dɈ��	�����$��FS�SOS��4h �6�zN5�%t"K"F2!d+���UsbC�e�Rb@�Mx�m��I�hфI���t�i n}�N�k�+�[���_W\τ��c�z���D��?���[����u�t6�|�v�]G�[��Z�����<{��$R����ͭ]x��(ؘ'~!�FS��W;�孕��qi����ɾ*�S�a����1�e�����+�&{]�|10`g�9���8�Л��e��	t�O�]�����Bms0�zѼ���rG9��W��єĩ��a�3�0�6���뾂��ɜ]�7z�.�u�w^
^�M�b�xuxbd�+�4�LM��i�Y�w�ޭ/yTR�n�j�$�"��I�48�EC:q���)�J�N�\��j0���$R�Ƀ�U4�E�cn�-�|j(�d�c�o<��{nf�)�;��՗����Cc��m��P���ptм��r�I�D�D�d:��r9�V���U�dM���#c1e0tBi#���3#X��(^��(F��\X�0����
o���Л��l��$9�����琣�h�ڨ9��@��N�Q1N���e%�f�8G[�3x糙��bW�G!�^���Hk���wdP�T'�Z38��q�{7�ܘ�
Z�t�#��F�J��1 Y�K3J������(��7<q>�E,����$��.�Z�Y=ZGA�۠z5]�f�ɬ$3��������3e0�;:���jm���dT���	ո�ǹ^��\5�9�K���7�z=�i~��Bu���J_;WGM�nm���<r���dQ$�Qj�t�]%"�Ht�����q���i��	ϯd�D�V+�x�8�Ɏ8����fxY!����w���ev��7`kyM���
W��l��\���W�o�@#e �GW:�(,�Ɩ:$#��a���=(��]�X��,#�Ғ%���[g7$�~h������&�Y�0��{�O�Q�h�=m"���gG:��L�]���ܨ���z�fK�+�f��"�v<�!4./�O&�N�sQ�M^lM{UR��:z�JG�����j3�C7��ژ�1��K��J4/!j��L Y6�����Q�uNY`�J_8U
�ul�m����R%N�e?��*��j(d��qz�0N�5\��LI��g>��~:���e��Қ*��f��w$S�	8^Q