BZh91AY&SYI�� �_�Px���������P��Zu9��L�0�4� h���P  �@5=h��0 L��� 0BDS�OF��2z2��  @0`��`ѐ��&��RH`L����Q=2��2 ��6�%t��F1#4!^�諵J����4*LAa"(S_�}�ۇM�CB�3�V�� '���׷�o��oc����3�3�ڪe��u���	��I(F����T��c�SF�%��0�j�*�X�f%�#���w��/Ա�zL%X��)��Õ��26Mծ�މ&f�K�&&��rIO�X��R���n6�m�9����p�$4��kwӬ9��2Y�fV��`��-�X�tR�k}�Ǡ��&�BHp��X3D�kHN0�j��S�j`Y!޸�
̴ˇe4�Z�g�&���&0�T��2�T[M����
��Ua*���M͝��`b�$���4h"PX`��D�Z�kg
�S.C�Æn��ag�G
��ڴqQ�f ��,cc��m�4�r��aߤ��d�RC���*Q%���1��#rF���@���"�*�QkH�dep!l�PP0�fغ��k;]3="~�/+�p���w,0��Z��,�&�mѪ���p�3�
h	��|w�R �a}�`.0Ds�ȣ����{Բ�Lv�z�G�p��흿��oa�L�E$��cY��^��R��R��m�M�t��#���L��@�I=)�ϖ	N����F��71=]Բ�k/�IZ�.��a�S5H�㭡�K7Rт�{p2�����p�(j`k6�Xc�S�N��-QW)��6L�idT�[k	����eدP�V���+��/K.�='��a�d��:�YaVnZyWG�����fݽz�v1Q��¢�F�ʸ(SNA��!/��	��ƺE(��ŋh�����1�Ύx��5T�n=	��h���-Q�;�٭����CZ�SkCݷ-Sl�gPjҠ�w�X�����H�d�7�b;B����S-/�Ѱwo�[�v�qp�j}:����>w���V��BŇW��v��MO=��6�%0�qp2]$W�j�Q�R���t���/w����/+��O����b����iR�*K�]��dj�m�����Jeh�A�8��̛�da/��<1h\�ֳ2���Щhmbp�re�q�J�Ņڬ�Y��r��vԋ�>u�c������>.c=y�ٜ�C"j�,��c��MT�8GH�D+Ah��'0{��ܑN$z� 