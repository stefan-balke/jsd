BZh91AY&SY��vY _�Px���������P>u�77:� xJM�L�I��F@��� �%4!����@4  h  �I	=@M��   sbh0�2d��`�i���!�H�)�&�Ƒ��S5=@ ��=4M���℈H�"���H��R�Z
`�&���o�b�B��0���ԛibr�OwN�\ܜ�v�����]&H�-�.vs�Y�O?TQ͌z�֤�����..0�W̘���N��挲>�C��[|��F�+�1��V�2 5�If�|�p����=�3��P:�4��v�˨<=����͜u
oW1:$ґ�s.&'*}�����[U��!�x0�,A�28�
p-�����/�t`�TFc ���eEf���b��u�қHiC_.N'HE���//a�@�}a%��՗g�ɮ[-�W�m��i[�7S�n���m��z�~�֘���NY$*��\��X8>+,�P���Ģ�ěiVQ��Dk��"4�roM����$G���]���thݬɘ/L��NZJ��0�<K��^�O���+b=�&G)A<��ʹ�����L=IZ����9����ck�?Hm�\�B����Gq�.�L;�����^�E���m�/�Ԩ������P\`609W�D)��`�v��s�f[l{�
����u�5K	�����1j�e̚71(9�L�)XR��\�p3ρc:��BCIƒ�6���? 4��)�0.5*
������|i�	�� �]������pd��L��k�6�M:	j���d�"�B�
Q�kB���@�	��������$D��v��H*J�%> ���`
��a���s�%�	�v��ra��Rr�Q!f 	�HPb��A������TAPZ�3�
s(T�$� �*��� "�m���j��W ^�2��ߥ"C�����&�@@�Pc��Q������0���B{�Ά� ���i	�f�*�Ǩ�/.⻦�@��s@�ۆHc(�^,�#�0׎aV[��sH�N�5'u���5�`�56hZ섂���xT@�C���i��涓�A���00�+ʥ�H���d8��_#j��������
���]��BBF��d