BZh91AY&SY�8�� <_�Pxg���������P9�fV��P���z�A���4 ��A� ��1%�       %=DAOQ��6� Ѡ  @dɦ�L����0Fh� 	� D�52��=F�S�@i�OPh&�:P�
���`�B���_��Y$y���hD�&I���6�3�ƅ`fP���BB�@f���5oj�]�߼��T�/Ǥ�g�NZRQ?~���������ݨV�Z3�������4UT����_����;�aPa��کi,F�L�4�Y�R�IA�싮����<�@�����BU3y����j`00)G<�NW�>��P8�M0c�o��}~��~�$�$��pQjQ��
;��<B��Ib$��Y�$t�v;o�k<d �<�KpL��#bg39
K5�N,��E��G&��Z�8Wh/��r��b� �U�1A��1T��$ڮ��L��K��I�J
U���+��Z�����8�T�ũ)H��f%l����,�T�jHgzR�C�P��-FS43����e���/$JE����/�0��!2�3l�d��<�(����I��:ݐ䨎]�Y�(�o=�&���U��^�9�]X�L()�E0%$I/2�UR�`��f�K�j�Έ���E��jHF"��)����)�6�p�)�>�O�a�d�gP������҆_ǜ�h�MA���~>���<�� �d�M-R�P�Jmi3��Ű�u�Ƃ%�(�>%�8=��J�C�� 1W�5a�SX2V@|�vD�¿F�IUH�I@�H��ST!����u�L��L�l*���k�OEU��3TX�������9f���E	t���)��s����0j��aJ�G{:�[:�yuL��BCI8�U*l~A�@d~m����LP%����S,�	tH5�[��$n����q�R�$1(`r��I�T�q�8�,k���֡�]����jV$��Ul���-��ѡ��]��#��������!�%�p�a���3HV�S���(���@:4� ��bdACI{H�D��9�p�s*M�P�ʉ(�"3��+�О���G0�,|Ѥ����
���8<�'0�ZN��6	��:�@X�~�4	4ut���	�Lݒ�X����+��3�Ӛs��ƅG���n�Fk��8��$[ ေ8]"��Rw��P�|�A�3��� �P8Q+�\H-a�q)-���J@e/b�&�y����dmi0OI�/`m�cj��KL��\�6�'K]��!��0�^�K��rE8P��8��