BZh91AY&SYaM�j _�Px���������Pt�� �� JMI�M6�zz��� 2  h5S�<)���4   h  �2�� �     �	���dɓ#	�i�F& �"@��I�)�MOi�<�d 3=&$�p� HT@���~�����hR
hL�^g�m����B�2�Pl��-��+O4��wB��nU�}��V�d��k���3�U�E��scnS�:M��de�=|�5�*2čC�#�0O�Ք�E ����<g�#R�z^
�s�T%d�����w����P8�4��ܾ�!���\.X��n�Li���d��j���%4<B��Ґ=	��ҧ$iC��	�n�.���}n���,,K�K]'
�X��ٗ��
uUX2j�N
Z�Pfd������$������1$��,�4D�!@!	K$�P"!���/l��piXM����DӢ�*h�������X����*Q$�I�Ɗq�$EKXHHC]8�6�4�,�dߧ�W�.��8)$������y��EY����d�m5�1�JxK\'�|)_���Q�KT�[gX:B;M���_��{C�X`4'����~��QL=`�\�Z��|�"���2�R^��r�2f��@�����y�Lm�d32���� �-�����[b_]M^��z�4Р͐��nj�e��H�"`�JH�gEqC��|KU��cm��q�C�0�W�}Gxۆ��30<�E �.Ӹ=��3ψ���a���$tU]5��� Ψh�������B���`.ju�d��t8z	n)��AA\��C)k[}����0A�L�gB�C�l3�`q�%�*05,S��iV5K�PDa�h�� ���历�1{�TH�^�6��2���(�"1ّ��mBz���Lj=��Hb��g���	�TyXdq� ���b�F�&ฐ����`�~��\�DL��W�:N���vuA��D��d�0�bH���Z6���5�ߠU�W߁���,N�5'~
!T�D@�fhZ�A��o�k�$���RZaQ����.Ƒ���j9�M/���I�^�։5�
�)"��<wb��6�Z��c�~�����H�
)��@